library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

entity Control is
PORT
   (
      sys_clk_i:                IN   std_logic;
      inst  :                   IN   std_logic_vector (7 DOWNTO 0) := "00000000";
      step  :                   IN   std_logic_vector (2 DOWNTO 0) := "000";
      flags :                   IN   std_logic_vector (7 DOWNTO 0) := "00000000";
      q_CONTROL16:              OUT  std_logic_vector (31 DOWNTO 0);
      q_HALT:                   OUT  std_logic := '0';
      q_MEM_ADDR_IN:            OUT  std_logic := '0';
      q_RAM_IN:                 OUT  std_logic := '0';
      q_RAM_OUT:                OUT  std_logic := '0';
      q_INST_OUT:               OUT  std_logic := '0';
      q_INST_IN:                OUT  std_logic := '0';
      q_A_IN:                   OUT  std_logic := '0';
      q_A_OUT:                  OUT  std_logic := '0';
      q_SUM_OUT:                OUT  std_logic := '0';
      q_SUBTRACT:               OUT  std_logic := '0';
      q_X_IN:                   OUT  std_logic := '0';
      q_X_OUT:                  OUT  std_logic := '0';
      q_Y_IN:                   OUT  std_logic := '0';
      q_Y_OUT:                  OUT  std_logic := '0';
      q_I_IN:                   OUT  std_logic := '0';           
      q_I_OUT:                  OUT  std_logic := '0';
      q_OUTREG_IN:              OUT  std_logic := '0';
      q_COUNTER_ENABLE:         OUT  std_logic := '0';
      q_COUNTER_OUT:            OUT  std_logic := '0';
      q_JUMP:                   OUT  std_logic := '0';
      q_FI:                     OUT  std_logic := '0';
      q_CurrentADDR:            OUT  std_logic_vector (12 downto 0) := "0000000000000"
   );
end Control;

architecture Behavioral of Control is

TYPE mem IS ARRAY(0 TO 8191) OF std_logic_vector(31 DOWNTO 0);
SIGNAL rom_block : mem := (others=> (others=>'0'));
signal addr: integer := 0;

signal q_HALT_t                     : std_logic := '0';
signal q_MEM_ADDR_IN_t              : std_logic := '0';
signal q_RAM_IN_t                   : std_logic := '0';
signal q_RAM_OUT_t                  : std_logic := '0';
signal q_INST_OUT_t                 : std_logic := '0';
signal q_INST_IN_t                  : std_logic := '0';
signal q_A_IN_t                     : std_logic := '0';
signal q_A_OUT_t                    : std_logic := '0';
signal q_SUM_OUT_t                  : std_logic := '0';
signal q_SUBTRACT_t                 : std_logic := '0';
signal q_X_IN_t                     : std_logic := '0';
signal q_X_OUT_t                    : std_logic := '0';
signal q_Y_IN_t                     : std_logic := '0';
signal q_Y_OUT_t                    : std_logic := '0';
signal q_I_IN_t                     : std_logic := '0';
signal q_I_OUT_t                    : std_logic := '0';
signal q_OUTREG_IN_t                : std_logic := '0';
signal q_COUNTER_ENABLE_t           : std_logic := '0';
signal q_COUNTER_OUT_t              : std_logic := '0';
signal q_JUMP_t                     : std_logic := '0';
signal q_FI_t                       : std_logic := '0';

begin
   --"ROM" programming   --TO DO, allow dynamic programming instead of hardcoding this...
   -- IOUT / IIN / YOUT / YIN / XOUT / HLT / MEMADDRIN / RAMIN / RAMOUT / INSTOUT / INSTIN / AIN / AOUT / SUMOUT / SUBTRACT / XIN / OUTREGIN / COUNTEN (PC++) / COUNTOUT (PC) / JUMP(set PC) / FI
                                                                   --INST       STEP   CF,ZF   
    
    rom_block(0)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(9)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(10)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(11)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(12)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(13)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(14)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(15)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(16)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(17)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(18)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(19)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(20)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(21)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(22)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(23)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(24)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(25)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(26)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(27)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(28)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(29)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(30)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(31)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(32)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(33)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(34)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(35)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(36)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(37)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(38)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(39)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(40)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(41)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(42)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(43)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(44)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(45)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(46)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(47)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(48)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(49)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(50)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(51)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(52)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(53)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(54)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(55)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(56)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(57)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(58)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(59)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(60)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(61)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(62)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(63)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(64)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(65)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(66)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(67)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(68)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(69)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(70)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(71)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(72)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(73)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(74)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(75)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(76)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(77)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(78)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(79)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(80)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(81)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(82)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(83)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(84)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(85)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(86)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(87)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(88)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(89)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(90)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(91)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(92)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(93)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(94)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(95)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(96)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(97)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(98)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(99)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(100)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(101)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(102)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(103)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(104)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(105)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(106)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(107)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(108)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(109)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(110)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(111)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(112)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(113)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(114)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(115)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(116)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(117)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(118)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(119)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(120)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(121)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(122)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(123)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(124)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(125)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(126)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(127)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(128)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(129)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(130)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(131)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(132)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(133)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(134)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(135)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(136)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(137)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(138)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(139)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(140)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(141)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(142)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(143)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(144)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(145)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(146)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(147)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(148)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(149)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(150)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(151)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(152)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(153)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(154)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(155)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(156)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(157)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(158)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(159)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(160)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(161)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(162)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(163)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(164)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(165)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(166)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(167)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(168)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(169)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(170)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(171)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(172)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(173)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(174)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(175)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(176)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(177)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(178)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(179)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(180)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(181)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(182)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(183)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(184)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(185)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(186)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(187)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(188)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(189)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(190)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(191)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(192)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(193)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(194)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(195)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(196)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(197)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(198)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(199)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(200)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(201)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(202)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(203)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(204)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(205)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(206)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(207)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(208)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(209)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(210)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(211)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(212)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(213)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(214)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(215)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(216)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(217)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(218)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(219)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(220)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(221)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(222)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(223)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(224)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(225)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(226)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(227)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(228)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(229)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(230)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(231)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(232)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(233)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(234)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(235)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(236)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(237)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(238)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(239)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(240)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(241)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(242)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(243)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(244)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(245)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(246)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(247)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(248)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(249)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(250)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(251)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(252)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(253)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(254)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(255)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(256)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(257)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(258)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(259)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(260)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(261)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(262)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(263)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(264)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(265)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(266)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(267)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(268)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(269)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(270)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(271)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(272)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(273)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(274)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(275)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(276)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(277)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(278)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(279)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(280)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(281)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(282)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(283)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(284)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(285)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(286)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(287)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(288)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(289)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(290)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(291)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(292)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(293)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(294)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(295)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(296)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(297)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(298)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(299)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(300)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(301)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(302)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(303)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(304)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(305)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(306)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(307)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(308)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(309)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(310)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(311)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(312)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(313)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(314)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(315)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(316)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(317)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(318)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(319)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(320)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(321)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(322)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(323)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(324)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(325)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(326)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(327)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(328)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(329)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(330)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(331)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(332)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(333)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(334)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(335)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(336)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(337)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(338)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(339)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(340)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(341)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(342)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(343)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(344)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(345)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(346)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(347)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(348)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(349)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(350)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(351)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(352)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(353)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(354)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(355)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(356)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(357)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(358)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(359)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(360)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(361)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(362)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(363)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(364)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(365)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(366)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(367)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(368)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(369)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(370)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(371)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(372)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(373)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(374)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(375)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(376)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(377)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(378)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(379)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(380)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(381)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(382)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(383)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(384)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(385)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(386)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(387)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(388)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(389)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(390)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(391)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(392)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(393)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(394)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(395)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(396)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(397)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(398)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(399)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(400)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(401)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(402)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(403)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(404)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(405)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(406)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(407)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(408)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(409)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(410)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(411)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(412)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(413)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(414)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(415)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(416)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(417)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(418)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(419)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(420)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(421)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(422)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(423)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(424)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(425)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(426)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(427)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(428)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(429)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(430)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(431)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(432)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(433)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(434)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(435)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(436)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(437)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(438)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(439)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(440)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(441)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(442)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(443)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(444)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(445)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(446)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(447)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(448)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(449)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(450)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(451)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(452)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(453)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(454)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(455)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(456)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(457)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(458)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(459)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(460)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(461)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(462)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(463)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(464)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(465)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(466)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(467)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(468)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(469)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(470)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(471)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(472)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(473)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(474)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(475)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(476)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(477)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(478)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(479)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(480)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(481)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(482)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(483)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(484)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(485)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(486)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(487)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(488)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(489)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(490)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(491)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(492)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(493)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(494)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(495)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(496)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(497)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(498)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(499)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(500)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(501)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(502)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(503)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(504)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(505)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(506)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(507)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(508)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(509)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(510)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(511)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(512)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(513)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(514)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(515)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(516)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(517)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(518)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(519)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(520)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(521)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(522)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(523)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(524)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(525)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(526)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(527)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(528)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(529)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(530)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(531)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(532)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(533)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(534)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(535)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(536)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(537)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(538)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(539)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(540)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(541)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(542)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(543)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(544)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(545)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(546)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(547)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(548)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(549)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(550)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(551)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(552)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(553)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(554)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(555)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(556)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(557)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(558)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(559)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(560)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(561)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(562)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(563)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(564)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(565)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(566)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(567)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(568)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(569)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(570)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(571)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(572)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(573)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(574)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(575)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(576)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(577)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(578)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(579)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(580)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(581)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(582)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(583)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(584)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(585)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(586)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(587)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(588)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(589)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(590)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(591)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(592)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(593)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(594)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(595)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(596)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(597)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(598)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(599)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(600)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(601)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(602)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(603)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(604)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(605)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(606)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(607)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(608)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(609)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(610)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(611)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(612)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(613)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(614)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(615)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(616)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(617)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(618)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(619)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(620)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(621)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(622)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(623)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(624)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(625)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(626)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(627)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(628)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(629)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(630)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(631)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(632)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(633)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(634)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(635)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(636)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(637)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(638)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(639)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(640)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(641)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(642)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(643)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(644)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(645)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(646)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(647)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(648)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(649)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(650)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(651)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(652)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(653)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(654)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(655)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(656)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(657)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(658)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(659)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(660)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(661)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(662)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(663)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(664)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(665)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(666)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(667)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(668)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(669)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(670)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(671)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(672)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(673)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(674)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(675)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(676)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(677)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(678)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(679)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(680)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(681)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(682)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(683)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(684)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(685)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(686)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(687)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(688)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(689)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(690)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(691)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(692)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(693)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(694)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(695)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(696)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(697)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(698)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(699)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(700)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(701)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(702)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(703)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(704)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(705)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(706)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(707)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(708)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(709)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(710)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(711)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(712)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(713)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(714)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(715)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(716)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(717)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(718)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(719)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(720)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(721)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(722)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(723)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(724)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(725)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(726)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(727)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(728)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(729)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(730)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(731)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(732)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(733)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(734)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(735)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(736)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(737)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(738)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(739)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(740)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(741)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(742)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(743)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(744)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(745)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(746)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(747)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(748)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(749)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(750)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(751)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(752)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(753)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(754)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(755)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(756)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(757)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(758)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(759)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(760)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(761)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(762)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(763)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(764)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(765)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(766)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(767)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(768)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(769)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(770)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(771)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(772)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(773)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(774)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(775)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(776)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(777)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(778)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(779)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(780)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(781)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(782)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(783)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(784)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(785)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(786)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(787)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(788)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(789)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(790)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(791)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(792)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(793)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(794)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(795)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(796)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(797)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(798)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(799)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(800)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(801)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(802)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(803)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(804)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(805)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(806)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(807)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(808)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(809)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(810)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(811)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(812)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(813)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(814)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(815)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(816)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(817)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(818)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(819)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(820)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(821)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(822)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(823)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(824)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(825)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(826)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(827)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(828)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(829)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(830)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(831)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(832)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(833)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(834)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(835)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(836)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(837)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(838)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(839)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(840)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(841)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(842)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(843)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(844)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(845)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(846)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(847)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(848)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(849)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(850)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(851)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(852)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(853)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(854)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(855)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(856)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(857)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(858)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(859)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(860)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(861)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(862)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(863)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(864)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(865)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(866)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(867)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(868)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(869)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(870)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(871)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(872)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(873)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(874)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(875)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(876)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(877)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(878)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(879)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(880)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(881)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(882)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(883)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(884)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(885)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(886)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(887)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(888)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(889)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(890)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(891)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(892)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(893)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(894)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(895)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(896)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(897)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(898)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(899)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(900)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(901)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(902)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(903)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(904)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(905)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(906)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(907)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(908)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(909)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(910)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(911)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(912)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(913)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(914)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(915)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(916)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(917)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(918)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(919)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(920)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(921)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(922)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(923)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(924)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(925)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(926)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(927)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(928)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(929)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(930)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(931)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(932)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(933)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(934)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(935)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(936)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(937)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(938)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(939)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(940)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(941)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(942)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(943)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(944)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(945)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(946)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(947)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(948)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(949)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(950)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(951)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(952)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(953)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(954)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(955)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(956)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(957)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(958)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(959)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(960)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(961)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(962)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(963)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(964)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(965)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(966)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(967)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(968)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(969)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(970)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(971)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(972)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(973)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(974)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(975)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(976)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(977)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(978)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(979)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(980)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(981)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(982)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(983)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(984)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(985)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(986)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(987)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(988)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(989)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(990)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(991)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(992)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(993)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(994)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(995)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(996)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(997)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(998)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(999)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1000)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1001)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1002)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1003)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1004)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1005)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1006)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1007)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1008)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1009)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1010)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1011)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1012)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1013)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1014)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1015)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1016)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1017)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1018)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1019)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1020)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1021)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1022)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1023)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1024)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1025)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1026)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1027)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1028)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1029)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1030)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1031)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1032)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1033)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1034)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1035)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1036)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1037)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1038)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1039)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1040)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1041)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1042)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1043)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1044)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1045)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1046)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1047)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1048)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1049)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1050)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1051)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1052)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1053)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1054)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1055)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1056)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1057)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1058)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1059)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1060)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1061)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1062)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1063)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1064)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1065)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1066)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1067)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1068)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1069)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1070)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1071)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1072)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1073)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1074)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1075)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1076)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1077)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1078)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1079)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1080)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1081)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1082)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1083)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1084)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1085)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1086)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1087)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1088)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1089)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1090)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1091)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1092)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1093)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1094)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1095)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1096)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1097)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1098)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1099)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1100)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1101)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1102)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1103)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1104)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1105)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1106)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1107)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1108)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1109)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1110)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1111)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1112)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1113)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1114)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1115)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1116)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1117)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1118)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1119)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1120)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1121)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1122)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1123)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1124)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1125)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1126)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1127)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1128)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1129)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1130)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1131)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1132)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1133)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1134)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1135)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1136)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1137)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1138)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1139)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1140)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1141)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1142)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1143)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1144)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1145)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1146)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1147)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1148)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1149)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1150)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1151)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1152)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1153)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1154)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1155)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1156)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1157)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1158)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1159)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1160)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1161)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1162)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1163)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1164)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1165)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1166)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1167)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1168)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1169)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1170)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1171)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1172)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1173)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1174)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1175)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1176)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1177)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1178)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1179)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1180)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1181)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1182)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1183)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1184)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1185)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1186)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1187)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1188)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1189)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1190)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1191)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1192)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1193)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1194)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1195)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1196)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1197)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1198)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1199)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1200)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1201)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1202)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1203)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1204)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1205)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1206)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1207)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1208)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1209)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1210)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1211)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1212)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1213)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1214)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1215)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1216)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1217)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1218)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1219)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1220)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1221)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1222)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1223)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1224)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1225)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1226)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1227)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1228)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1229)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1230)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1231)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1232)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1233)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1234)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1235)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1236)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1237)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1238)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1239)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1240)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1241)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1242)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1243)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1244)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1245)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1246)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1247)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1248)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1249)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1250)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1251)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1252)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1253)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1254)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1255)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1256)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1257)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1258)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1259)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1260)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1261)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1262)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1263)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1264)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1265)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1266)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1267)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1268)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1269)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1270)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1271)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1272)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1273)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1274)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1275)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1276)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1277)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1278)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1279)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1280)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1281)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1282)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1283)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1284)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1285)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1286)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1287)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1288)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1289)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1290)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1291)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1292)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1293)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1294)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1295)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1296)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1297)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1298)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1299)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1300)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1301)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1302)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1303)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1304)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1305)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1306)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1307)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1308)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1309)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1310)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1311)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1312)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1313)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1314)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1315)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1316)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1317)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1318)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1319)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1320)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1321)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1322)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1323)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1324)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1325)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1326)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1327)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1328)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1329)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1330)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1331)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1332)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1333)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1334)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1335)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1336)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1337)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1338)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1339)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1340)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1341)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1342)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1343)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1344)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1345)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1346)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1347)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1348)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1349)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1350)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1351)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1352)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1353)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1354)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1355)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1356)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1357)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1358)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1359)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1360)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1361)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1362)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1363)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1364)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1365)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1366)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1367)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1368)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1369)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1370)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1371)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1372)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1373)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1374)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1375)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1376)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1377)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1378)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1379)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1380)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1381)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1382)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1383)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1384)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1385)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1386)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1387)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1388)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1389)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1390)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1391)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1392)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1393)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1394)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1395)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1396)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1397)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1398)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1399)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1400)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1401)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1402)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1403)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1404)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1405)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1406)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1407)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1408)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1409)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1410)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1411)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1412)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1413)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1414)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1415)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1416)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1417)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1418)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1419)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1420)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1421)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1422)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1423)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1424)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1425)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1426)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1427)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1428)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1429)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1430)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1431)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1432)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1433)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1434)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1435)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1436)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1437)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1438)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1439)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1440)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1441)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1442)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1443)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1444)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1445)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1446)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1447)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1448)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1449)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1450)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1451)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1452)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1453)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1454)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1455)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1456)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1457)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1458)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1459)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1460)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1461)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1462)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1463)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1464)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1465)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1466)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1467)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1468)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1469)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1470)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1471)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1472)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1473)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1474)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1475)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1476)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1477)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1478)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1479)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1480)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1481)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1482)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1483)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1484)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1485)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1486)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1487)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1488)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1489)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1490)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1491)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1492)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1493)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1494)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1495)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1496)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1497)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1498)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1499)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1500)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1501)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1502)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1503)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1504)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1505)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1506)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1507)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1508)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1509)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1510)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1511)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1512)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1513)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1514)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1515)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1516)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1517)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1518)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1519)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1520)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1521)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1522)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1523)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1524)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1525)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1526)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1527)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1528)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1529)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1530)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1531)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1532)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1533)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1534)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1535)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1536)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1537)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1538)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1539)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1540)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1541)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1542)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1543)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1544)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1545)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1546)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1547)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1548)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1549)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1550)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1551)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1552)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1553)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1554)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1555)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1556)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1557)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1558)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1559)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1560)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1561)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1562)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1563)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1564)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1565)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1566)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1567)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1568)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1569)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1570)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1571)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1572)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1573)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1574)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1575)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1576)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1577)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1578)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1579)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1580)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1581)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1582)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1583)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1584)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1585)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1586)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1587)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1588)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1589)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1590)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1591)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1592)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1593)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1594)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1595)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1596)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1597)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1598)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1599)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1600)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1601)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1602)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1603)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1604)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1605)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1606)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1607)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1608)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1609)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1610)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1611)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1612)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1613)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1614)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1615)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1616)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1617)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1618)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1619)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1620)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1621)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1622)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1623)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1624)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1625)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1626)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1627)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1628)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1629)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1630)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1631)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1632)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1633)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1634)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1635)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1636)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1637)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1638)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1639)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1640)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1641)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1642)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1643)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1644)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1645)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1646)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1647)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1648)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1649)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1650)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1651)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1652)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1653)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1654)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1655)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1656)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1657)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1658)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1659)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1660)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1661)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1662)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1663)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1664)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1665)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1666)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1667)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1668)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1669)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1670)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1671)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1672)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1673)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1674)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1675)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1676)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1677)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1678)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1679)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1680)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1681)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1682)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1683)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1684)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1685)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1686)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1687)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1688)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1689)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1690)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1691)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1692)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1693)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1694)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1695)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1696)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1697)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1698)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1699)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1700)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1701)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1702)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1703)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1704)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1705)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1706)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1707)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1708)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1709)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1710)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1711)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1712)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1713)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1714)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1715)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1716)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1717)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1718)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1719)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1720)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1721)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1722)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1723)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1724)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1725)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1726)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1727)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1728)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1729)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1730)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1731)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1732)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1733)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1734)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1735)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1736)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1737)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1738)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1739)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1740)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1741)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1742)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1743)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1744)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1745)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1746)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1747)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1748)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1749)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1750)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1751)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1752)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1753)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1754)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1755)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1756)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1757)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1758)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1759)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1760)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1761)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1762)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1763)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1764)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1765)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1766)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1767)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1768)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1769)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1770)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1771)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1772)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1773)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1774)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1775)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1776)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1777)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1778)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1779)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1780)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1781)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1782)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1783)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1784)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1785)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1786)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1787)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1788)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1789)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1790)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1791)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1792)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1793)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1794)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1795)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1796)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1797)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1798)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1799)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1800)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1801)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1802)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1803)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1804)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1805)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1806)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1807)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1808)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1809)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1810)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1811)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1812)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1813)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1814)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1815)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1816)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1817)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1818)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1819)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1820)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1821)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1822)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1823)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1824)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1825)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1826)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1827)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1828)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1829)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1830)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1831)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1832)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1833)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1834)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1835)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1836)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1837)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1838)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1839)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1840)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1841)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1842)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1843)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1844)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1845)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1846)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1847)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1848)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1849)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1850)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1851)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1852)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1853)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1854)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1855)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1856)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1857)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1858)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1859)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1860)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1861)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1862)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1863)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1864)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1865)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1866)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1867)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1868)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1869)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1870)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1871)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1872)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1873)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1874)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1875)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1876)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1877)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1878)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1879)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1880)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1881)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1882)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1883)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1884)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1885)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1886)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1887)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1888)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1889)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1890)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1891)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1892)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1893)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1894)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1895)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1896)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1897)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1898)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1899)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1900)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1901)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1902)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1903)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1904)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1905)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1906)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1907)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1908)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1909)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1910)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1911)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1912)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1913)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1914)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1915)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1916)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1917)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1918)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1919)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1920)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1921)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1922)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1923)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1924)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1925)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1926)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1927)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1928)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1929)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1930)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1931)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1932)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1933)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1934)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1935)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1936)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1937)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1938)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1939)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(1940)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1941)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1942)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1943)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(1944)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1945)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1946)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1947)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(1948)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1949)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1950)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1951)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(1952)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1953)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1954)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1955)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(1956)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1957)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1958)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1959)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(1960)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1961)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1962)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1963)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(1964)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1965)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1966)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1967)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(1968)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1969)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1970)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1971)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(1972)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1973)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1974)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1975)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(1976)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1977)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1978)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1979)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(1980)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1981)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1982)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1983)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(1984)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1985)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1986)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1987)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(1988)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1989)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1990)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1991)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(1992)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1993)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1994)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1995)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(1996)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1997)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1998)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(1999)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2000)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2001)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2002)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2003)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2004)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2005)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2006)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2007)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2008)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2009)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2010)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2011)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2012)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2013)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2014)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2015)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2016)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2017)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2018)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2019)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2020)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2021)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2022)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2023)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2024)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2025)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2026)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2027)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2028)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2029)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2030)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2031)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2032)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2033)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2034)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2035)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2036)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2037)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2038)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2039)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2040)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2041)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2042)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2043)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2044)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2045)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2046)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2047)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2048)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2049)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2050)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2051)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2052)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2053)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2054)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2055)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2056)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2057)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2058)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2059)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2060)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2061)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2062)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2063)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2064)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2065)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2066)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2067)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2068)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2069)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2070)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2071)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2072)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2073)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2074)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2075)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2076)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2077)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2078)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2079)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2080)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2081)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2082)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2083)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2084)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2085)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2086)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2087)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2088)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2089)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2090)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2091)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2092)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2093)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2094)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2095)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2096)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2097)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2098)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2099)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2100)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2101)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2102)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2103)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2104)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2105)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2106)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2107)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2108)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2109)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2110)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2111)   <="00000000000000000000000000000000";    --TBD2:7
    
    --HLT / MEMADDRIN / RAMIN / RAMOUT / INSTOUT / INSTIN / AIN / AOUT / SUMOUT / SUBTRACT / BIN / OUTREGIN / COUNTEN (PC++) / COUNTOUT (PC) / JUMP(set PC) / FI
    --JMPA (42)
    rom_block(2112)   <="00000000000000000100000000000100";    --JMPA:0 (WDM reserved)
    rom_block(2113)   <="00000000000000000100000000000100";    --JMPA:0
    rom_block(2114)   <="00000000000000000100000000000100";    --JMPA:0
    rom_block(2115)   <="00000000000000000100000000000100";    --JMPA:0
    rom_block(2116)   <="00000000000000000001010000001000";    --JMPA:1
    rom_block(2117)   <="00000000000000000001010000001000";    --JMPA:1
    rom_block(2118)   <="00000000000000000001010000001000";    --JMPA:1
    rom_block(2119)   <="00000000000000000001010000001000";    --JMPA:1
    rom_block(2120)   <="00000000000000000000000100001010";    --JMPA:2  --** calling JMP twice, as the Vivado IP for binary counter load applies to the next clock rise. CE must also be high during the read of new values.
    rom_block(2121)   <="00000000000000000000000100001010";    --JMPA:2
    rom_block(2122)   <="00000000000000000000000100001010";    --JMPA:2
    rom_block(2123)   <="00000000000000000000000100001010";    --JMPA:2
    rom_block(2124)   <="00000000000000000000000100001010";    --JMPA:3
    rom_block(2125)   <="00000000000000000000000100001010";    --JMPA:3
    rom_block(2126)   <="00000000000000000000000100001010";    --JMPA:3
    rom_block(2127)   <="00000000000000000000000100001010";    --JMPA:3
    rom_block(2128)   <="00000000000000000000000000000000";    --JMPA:4
    rom_block(2129)   <="00000000000000000000000000000000";    --JMPA:4
    rom_block(2130)   <="00000000000000000000000000000000";    --JMPA:4
    rom_block(2131)   <="00000000000000000000000000000000";    --JMPA:4
    rom_block(2132)   <="00000000000000000000000000000000";    --JMPA:5
    rom_block(2133)   <="00000000000000000000000000000000";    --JMPA:5
    rom_block(2134)   <="00000000000000000000000000000000";    --JMPA:5
    rom_block(2135)   <="00000000000000000000000000000000";    --JMPA:5
    rom_block(2136)   <="00000000000000000000000000000000";    --JMPA:6
    rom_block(2137)   <="00000000000000000000000000000000";    --JMPA:6
    rom_block(2138)   <="00000000000000000000000000000000";    --JMPA:6
    rom_block(2139)   <="00000000000000000000000000000000";    --JMPA:6
    rom_block(2140)   <="00000000000000000000000000000000";    --JMPA:7
    rom_block(2141)   <="00000000000000000000000000000000";    --JMPA:7
    rom_block(2142)   <="00000000000000000000000000000000";    --JMPA:7
    rom_block(2143)   <="00000000000000000000000000000000";    --JMPA:7
    
    rom_block(2144)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2145)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2146)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2147)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2148)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2149)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2150)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2151)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2152)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2153)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2154)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2155)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2156)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2157)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2158)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2159)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2160)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2161)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2162)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2163)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2164)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2165)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2166)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2167)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2168)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2169)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2170)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2171)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2172)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2173)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2174)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2175)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2176)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2177)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2178)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2179)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2180)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2181)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2182)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2183)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2184)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2185)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2186)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2187)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2188)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2189)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2190)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2191)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2192)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2193)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2194)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2195)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2196)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2197)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2198)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2199)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2200)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2201)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2202)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2203)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2204)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2205)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2206)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2207)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2208)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2209)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2210)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2211)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2212)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2213)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2214)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2215)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2216)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2217)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2218)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2219)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2220)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2221)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2222)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2223)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2224)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2225)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2226)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2227)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2228)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2229)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2230)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2231)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2232)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2233)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2234)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2235)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2236)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2237)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2238)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2239)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2240)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2241)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2242)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2243)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2244)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2245)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2246)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2247)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2248)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2249)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2250)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2251)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2252)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2253)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2254)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2255)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2256)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2257)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2258)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2259)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2260)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2261)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2262)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2263)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2264)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2265)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2266)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2267)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2268)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2269)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2270)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2271)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2272)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2273)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2274)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2275)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2276)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2277)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2278)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2279)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2280)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2281)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2282)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2283)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2284)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2285)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2286)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2287)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2288)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2289)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2290)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2291)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2292)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2293)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2294)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2295)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2296)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2297)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2298)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2299)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2300)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2301)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2302)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2303)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2304)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2305)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2306)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2307)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2308)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2309)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2310)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2311)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2312)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2313)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2314)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2315)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2316)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2317)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2318)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2319)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2320)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2321)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2322)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2323)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2324)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2325)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2326)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2327)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2328)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2329)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2330)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2331)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2332)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2333)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2334)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2335)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2336)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2337)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2338)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2339)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2340)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2341)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2342)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2343)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2344)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2345)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2346)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2347)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2348)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2349)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2350)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2351)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2352)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2353)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2354)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2355)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2356)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2357)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2358)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2359)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2360)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2361)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2362)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2363)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2364)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2365)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2366)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2367)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2368)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2369)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2370)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2371)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2372)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2373)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2374)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2375)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2376)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2377)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2378)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2379)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2380)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2381)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2382)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2383)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2384)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2385)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2386)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2387)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2388)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2389)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2390)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2391)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2392)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2393)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2394)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2395)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2396)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2397)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2398)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2399)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2400)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2401)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2402)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2403)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2404)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2405)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2406)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2407)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2408)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2409)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2410)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2411)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2412)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2413)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2414)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2415)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2416)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2417)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2418)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2419)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2420)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2421)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2422)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2423)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2424)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2425)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2426)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2427)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2428)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2429)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2430)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2431)   <="00000000000000000000000000000000";    --TBD2:7

	-- xx/xx/xx/xx/xx/xx/xx/xx
    -- xx/xx/xx/ IOUT / IIN / YOUT / YIN / XOUT 
    -- HLT / MEMADDRIN / RAMIN / RAMOUT / INSTOUT / INSTIN / AIN / AOUT 
    -- SUMOUT / SUBTRACT / XIN / OUTREGIN / COUNTEN (PC++) / COUNTOUT (PC) / JUMP(set PC) / FI   
        
    --JMP (4C)
    rom_block(2432)   <="00000000000000000100000000000100";    --JMP:0      01001100  000 00
    rom_block(2433)   <="00000000000000000100000000000100";    --JMP:0
    rom_block(2434)   <="00000000000000000100000000000100";    --JMP:0
    rom_block(2435)   <="00000000000000000100000000000100";    --JMP:0
    rom_block(2436)   <="00000000000000000001010000001000";    --JMP:1
    rom_block(2437)   <="00000000000000000001010000001000";    --JMP:1
    rom_block(2438)   <="00000000000000000001010000001000";    --JMP:1
    rom_block(2439)   <="00000000000000000001010000001000";    --JMP:1
    rom_block(2440)   <=B"0000000000000000_01000000_00000100";    --JMP:2
    rom_block(2441)   <=B"0000000000000000_01000000_00000100";    --JMP:2
    rom_block(2442)   <=B"0000000000000000_01000000_00000100";    --JMP:2
    rom_block(2443)   <=B"0000000000000000_01000000_00000100";    --JMP:2
    rom_block(2444)   <=B"00000000_00001000_00010000_00001000";    --JMP:3
    rom_block(2445)   <=B"00000000_00001000_00010000_00001000";    --JMP:3
    rom_block(2446)   <=B"00000000_00001000_00010000_00001000";    --JMP:3
    rom_block(2447)   <=B"00000000_00001000_00010000_00001000";    --JMP:3
    rom_block(2448)   <=B"00000000_00010000_00000000_00001010";    --JMP:4  --** calling JMP twice, as the Vivado IP for binary counter load applies to the next clock rise. CE must also be high during the read of new values.
    rom_block(2449)   <=B"00000000_00010000_00000000_00001010";    --JMP:4
    rom_block(2450)   <=B"00000000_00010000_00000000_00001010";    --JMP:4
    rom_block(2451)   <=B"00000000_00010000_00000000_00001010";    --JMP:4
    rom_block(2452)   <=B"00000000_00010000_00000000_00001010";    --JMP:5
    rom_block(2453)   <=B"00000000_00010000_00000000_00001010";    --JMP:5
    rom_block(2454)   <=B"00000000_00010000_00000000_00001010";    --JMP:5
    rom_block(2455)   <=B"00000000_00010000_00000000_00001010";    --JMP:5
    rom_block(2456)   <="00000000000000000000000000000000";    --JMP:6
    rom_block(2457)   <="00000000000000000000000000000000";    --JMP:6
    rom_block(2458)   <="00000000000000000000000000000000";    --JMP:6
    rom_block(2459)   <="00000000000000000000000000000000";    --JMP:6
    rom_block(2460)   <="00000000000000000000000000000000";    --JMP:7
    rom_block(2461)   <="00000000000000000000000000000000";    --JMP:7
    rom_block(2462)   <="00000000000000000000000000000000";    --JMP:7
    rom_block(2463)   <="00000000000000000000000000000000";    --JMP:7
    rom_block(2464)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2465)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2466)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2467)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2468)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2469)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2470)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2471)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2472)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2473)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2474)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2475)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2476)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2477)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2478)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2479)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2480)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2481)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2482)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2483)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2484)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2485)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2486)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2487)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2488)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2489)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2490)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2491)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2492)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2493)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2494)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2495)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2496)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2497)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2498)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2499)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2500)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2501)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2502)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2503)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2504)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2505)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2506)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2507)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2508)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2509)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2510)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2511)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2512)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2513)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2514)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2515)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2516)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2517)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2518)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2519)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2520)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2521)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2522)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2523)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2524)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2525)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2526)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2527)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2528)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2529)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2530)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2531)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2532)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2533)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2534)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2535)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2536)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2537)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2538)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2539)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2540)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2541)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2542)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2543)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2544)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2545)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2546)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2547)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2548)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2549)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2550)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2551)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2552)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2553)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2554)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2555)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2556)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2557)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2558)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2559)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2560)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2561)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2562)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2563)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2564)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2565)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2566)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2567)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2568)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2569)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2570)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2571)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2572)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2573)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2574)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2575)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2576)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2577)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2578)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2579)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2580)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2581)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2582)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2583)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2584)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2585)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2586)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2587)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2588)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2589)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2590)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2591)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2592)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2593)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2594)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2595)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2596)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2597)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2598)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2599)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2600)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2601)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2602)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2603)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2604)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2605)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2606)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2607)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2608)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2609)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2610)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2611)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2612)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2613)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2614)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2615)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2616)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2617)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2618)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2619)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2620)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2621)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2622)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2623)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2624)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2625)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2626)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2627)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2628)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2629)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2630)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2631)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2632)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2633)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2634)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2635)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2636)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2637)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2638)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2639)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2640)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2641)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2642)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2643)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2644)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2645)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2646)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2647)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2648)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2649)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2650)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2651)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2652)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2653)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2654)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2655)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2656)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2657)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2658)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2659)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2660)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2661)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2662)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2663)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2664)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2665)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2666)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2667)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2668)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2669)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2670)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2671)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2672)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2673)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2674)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2675)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2676)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2677)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2678)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2679)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2680)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2681)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2682)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2683)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2684)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2685)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2686)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2687)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2688)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2689)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2690)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2691)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2692)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2693)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2694)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2695)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2696)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2697)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2698)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2699)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2700)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2701)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2702)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2703)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2704)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2705)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2706)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2707)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2708)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2709)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2710)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2711)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2712)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2713)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2714)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2715)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2716)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2717)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2718)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2719)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2720)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2721)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2722)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2723)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2724)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2725)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2726)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2727)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2728)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2729)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2730)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2731)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2732)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2733)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2734)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2735)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2736)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2737)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2738)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2739)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2740)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2741)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2742)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2743)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2744)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2745)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2746)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2747)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2748)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2749)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2750)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2751)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2752)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2753)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2754)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2755)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2756)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2757)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2758)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2759)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2760)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2761)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2762)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2763)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2764)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2765)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2766)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2767)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2768)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2769)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2770)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2771)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2772)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2773)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2774)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2775)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2776)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2777)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2778)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2779)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2780)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2781)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2782)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2783)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2784)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2785)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2786)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2787)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2788)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2789)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2790)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2791)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2792)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2793)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2794)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2795)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2796)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2797)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2798)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2799)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2800)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2801)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2802)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2803)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2804)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2805)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2806)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2807)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2808)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2809)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2810)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2811)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2812)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2813)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2814)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2815)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2816)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2817)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2818)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2819)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2820)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2821)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2822)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2823)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2824)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2825)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2826)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2827)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2828)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2829)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2830)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2831)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2832)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2833)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2834)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2835)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2836)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2837)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2838)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2839)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2840)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2841)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2842)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2843)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2844)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2845)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2846)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2847)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2848)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2849)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2850)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2851)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2852)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2853)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2854)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2855)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2856)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2857)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2858)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2859)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2860)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2861)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2862)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2863)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2864)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2865)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2866)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2867)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2868)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2869)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2870)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2871)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2872)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2873)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2874)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2875)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2876)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2877)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2878)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2879)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2880)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2881)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2882)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2883)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2884)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2885)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2886)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2887)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2888)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2889)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2890)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2891)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2892)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2893)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2894)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2895)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2896)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2897)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2898)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2899)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2900)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2901)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2902)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2903)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2904)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2905)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2906)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2907)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2908)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2909)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2910)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2911)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2912)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2913)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2914)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2915)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2916)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2917)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2918)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2919)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2920)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2921)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2922)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2923)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2924)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2925)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2926)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2927)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2928)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2929)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2930)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2931)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2932)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2933)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2934)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2935)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2936)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2937)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2938)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2939)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(2940)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2941)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2942)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2943)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(2944)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2945)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2946)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2947)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(2948)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2949)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2950)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2951)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(2952)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2953)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2954)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2955)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(2956)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2957)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2958)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2959)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(2960)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2961)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2962)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2963)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(2964)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2965)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2966)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2967)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(2968)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2969)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2970)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2971)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(2972)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2973)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2974)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2975)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(2976)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2977)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2978)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2979)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(2980)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2981)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2982)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2983)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(2984)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2985)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2986)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2987)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(2988)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2989)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2990)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2991)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(2992)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2993)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2994)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2995)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(2996)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2997)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2998)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(2999)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3000)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3001)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3002)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3003)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3004)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3005)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3006)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3007)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3008)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3009)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3010)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3011)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3012)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3013)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3014)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3015)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3016)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3017)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3018)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3019)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3020)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3021)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3022)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3023)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3024)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3025)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3026)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3027)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3028)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3029)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3030)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3031)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3032)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3033)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3034)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3035)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3036)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3037)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3038)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3039)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3040)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3041)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3042)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3043)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3044)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3045)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3046)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3047)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3048)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3049)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3050)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3051)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3052)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3053)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3054)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3055)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3056)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3057)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3058)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3059)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3060)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3061)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3062)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3063)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3064)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3065)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3066)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3067)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3068)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3069)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3070)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3071)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3072)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3073)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3074)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3075)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3076)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3077)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3078)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3079)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3080)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3081)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3082)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3083)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3084)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3085)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3086)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3087)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3088)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3089)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3090)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3091)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3092)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3093)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3094)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3095)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3096)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3097)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3098)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3099)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3100)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3101)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3102)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3103)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3104)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3105)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3106)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3107)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3108)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3109)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3110)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3111)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3112)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3113)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3114)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3115)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3116)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3117)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3118)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3119)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3120)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3121)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3122)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3123)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3124)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3125)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3126)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3127)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3128)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3129)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3130)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3131)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3132)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3133)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3134)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3135)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3136)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3137)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3138)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3139)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3140)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3141)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3142)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3143)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3144)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3145)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3146)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3147)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3148)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3149)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3150)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3151)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3152)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3153)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3154)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3155)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3156)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3157)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3158)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3159)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3160)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3161)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3162)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3163)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3164)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3165)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3166)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3167)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3168)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3169)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3170)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3171)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3172)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3173)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3174)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3175)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3176)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3177)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3178)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3179)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3180)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3181)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3182)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3183)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3184)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3185)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3186)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3187)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3188)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3189)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3190)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3191)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3192)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3193)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3194)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3195)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3196)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3197)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3198)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3199)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3200)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3201)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3202)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3203)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3204)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3205)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3206)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3207)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3208)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3209)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3210)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3211)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3212)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3213)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3214)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3215)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3216)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3217)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3218)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3219)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3220)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3221)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3222)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3223)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3224)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3225)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3226)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3227)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3228)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3229)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3230)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3231)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3232)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3233)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3234)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3235)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3236)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3237)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3238)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3239)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3240)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3241)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3242)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3243)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3244)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3245)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3246)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3247)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3248)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3249)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3250)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3251)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3252)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3253)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3254)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3255)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3256)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3257)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3258)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3259)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3260)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3261)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3262)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3263)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3264)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3265)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3266)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3267)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3268)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3269)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3270)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3271)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3272)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3273)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3274)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3275)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3276)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3277)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3278)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3279)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3280)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3281)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3282)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3283)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3284)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3285)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3286)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3287)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3288)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3289)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3290)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3291)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3292)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3293)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3294)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3295)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3296)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3297)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3298)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3299)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3300)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3301)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3302)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3303)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3304)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3305)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3306)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3307)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3308)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3309)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3310)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3311)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3312)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3313)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3314)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3315)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3316)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3317)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3318)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3319)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3320)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3321)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3322)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3323)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3324)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3325)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3326)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3327)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3328)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3329)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3330)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3331)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3332)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3333)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3334)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3335)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3336)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3337)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3338)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3339)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3340)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3341)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3342)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3343)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3344)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3345)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3346)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3347)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3348)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3349)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3350)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3351)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3352)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3353)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3354)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3355)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3356)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3357)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3358)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3359)   <="00000000000000000000000000000000";    --TBD:7
    
    -- xx/xx/xx/xx/xx/xx/xx/xx
    -- xx/xx/xx/ IOUT / IIN / YOUT / YIN / XOUT 
    -- HLT / MEMADDRIN / RAMIN / RAMOUT / INSTOUT / INSTIN / AIN / AOUT 
    -- SUMOUT / SUBTRACT / XIN / OUTREGIN / COUNTEN (PC++) / COUNTOUT (PC) / JUMP(set PC) / FI   
    
    --ADC Immed (69)
    rom_block(3360)   <="00000000000000000100000000000100";    --ADCI:0
    rom_block(3361)   <="00000000000000000100000000000100";    --ADCI:0
    rom_block(3362)   <="00000000000000000100000000000100";    --ADCI:0
    rom_block(3363)   <="00000000000000000100000000000100";    --ADCI:0
    rom_block(3364)   <="00000000000000000001010000001000";    --ADCI:1
    rom_block(3365)   <="00000000000000000001010000001000";    --ADCI:1
    rom_block(3366)   <="00000000000000000001010000001000";    --ADCI:1
    rom_block(3367)   <="00000000000000000001010000001000";    --ADCI:1
    rom_block(3368)   <=B"0000000000000000_0100000000000100";    --ADCI:2
    rom_block(3369)   <=B"0000000000000000_0100000000000100";    --ADCI:2
    rom_block(3370)   <=B"0000000000000000_0100000000000100";    --ADCI:2
    rom_block(3371)   <=B"0000000000000000_0100000000000100";    --ADCI:2
    rom_block(3372)   <=B"0000000000001000_0001000000001000";    --ADCI:3
    rom_block(3373)   <=B"0000000000001000_0001000000001000";    --ADCI:3
    rom_block(3374)   <=B"0000000000001000_0001000000001000";    --ADCI:3
    rom_block(3375)   <=B"0000000000001000_0001000000001000";    --ADCI:3
    rom_block(3376)   <=B"0000000000000000_00000010_10000001";    --ADCI:4
    rom_block(3377)   <=B"0000000000000000_00000010_10000001";    --ADCI:4
    rom_block(3378)   <=B"0000000000000000_00000010_10000001";    --ADCI:4
    rom_block(3379)   <=B"0000000000000000_00000010_10000001";    --ADCI:4
    rom_block(3380)   <="00000000000000000000000000000100";    --ADCI:5
    rom_block(3381)   <="00000000000000000000000000000100";    --ADCI:5
    rom_block(3382)   <="00000000000000000000000000000100";    --ADCI:5
    rom_block(3383)   <="00000000000000000000000000000100";    --ADCI:5
    rom_block(3384)   <="00000000000000000000000000000000";    --ADCI:6
    rom_block(3385)   <="00000000000000000000000000000000";    --ADCI:6
    rom_block(3386)   <="00000000000000000000000000000000";    --ADCI:6
    rom_block(3387)   <="00000000000000000000000000000000";    --ADCI:6
    rom_block(3388)   <="00000000000000000000000000000000";    --ADCI:7
    rom_block(3389)   <="00000000000000000000000000000000";    --ADCI:7
    rom_block(3390)   <="00000000000000000000000000000000";    --ADCI:7
    rom_block(3391)   <="00000000000000000000000000000000";    --ADCI:7
    
    rom_block(3392)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3393)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3394)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3395)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3396)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3397)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3398)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3399)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3400)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3401)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3402)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3403)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3404)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3405)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3406)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3407)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3408)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3409)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3410)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3411)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3412)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3413)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3414)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3415)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3416)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3417)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3418)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3419)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3420)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3421)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3422)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3423)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3424)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3425)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3426)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3427)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3428)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3429)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3430)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3431)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3432)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3433)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3434)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3435)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3436)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3437)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3438)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3439)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3440)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3441)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3442)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3443)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3444)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3445)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3446)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3447)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3448)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3449)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3450)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3451)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3452)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3453)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3454)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3455)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3456)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3457)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3458)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3459)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3460)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3461)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3462)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3463)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3464)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3465)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3466)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3467)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3468)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3469)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3470)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3471)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3472)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3473)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3474)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3475)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3476)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3477)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3478)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3479)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3480)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3481)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3482)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3483)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3484)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3485)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3486)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3487)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3488)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3489)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3490)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3491)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3492)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3493)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3494)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3495)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3496)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3497)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3498)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3499)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3500)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3501)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3502)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3503)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3504)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3505)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3506)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3507)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3508)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3509)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3510)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3511)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3512)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3513)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3514)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3515)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3516)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3517)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3518)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3519)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3520)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3521)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3522)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3523)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3524)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3525)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3526)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3527)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3528)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3529)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3530)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3531)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3532)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3533)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3534)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3535)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3536)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3537)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3538)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3539)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3540)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3541)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3542)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3543)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3544)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3545)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3546)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3547)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3548)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3549)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3550)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3551)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3552)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3553)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3554)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3555)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3556)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3557)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3558)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3559)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3560)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3561)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3562)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3563)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3564)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3565)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3566)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3567)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3568)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3569)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3570)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3571)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3572)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3573)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3574)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3575)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3576)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3577)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3578)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3579)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3580)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3581)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3582)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3583)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3584)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3585)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3586)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3587)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3588)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3589)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3590)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3591)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3592)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3593)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3594)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3595)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3596)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3597)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3598)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3599)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3600)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3601)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3602)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3603)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3604)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3605)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3606)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3607)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3608)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3609)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3610)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3611)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3612)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3613)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3614)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3615)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3616)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3617)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3618)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3619)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3620)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3621)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3622)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3623)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3624)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3625)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3626)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3627)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3628)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3629)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3630)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3631)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3632)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3633)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3634)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3635)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3636)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3637)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3638)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3639)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3640)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3641)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3642)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3643)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3644)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3645)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3646)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3647)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3648)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3649)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3650)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3651)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3652)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3653)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3654)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3655)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3656)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3657)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3658)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3659)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3660)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3661)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3662)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3663)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3664)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3665)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3666)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3667)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3668)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3669)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3670)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3671)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3672)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3673)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3674)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3675)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3676)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3677)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3678)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3679)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3680)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3681)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3682)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3683)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3684)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3685)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3686)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3687)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3688)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3689)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3690)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3691)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3692)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3693)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3694)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3695)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3696)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3697)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3698)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3699)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3700)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3701)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3702)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3703)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3704)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3705)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3706)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3707)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3708)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3709)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3710)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3711)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3712)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3713)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3714)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3715)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3716)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3717)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3718)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3719)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3720)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3721)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3722)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3723)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3724)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3725)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3726)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3727)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3728)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3729)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3730)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3731)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3732)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3733)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3734)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3735)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3736)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3737)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3738)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3739)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3740)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3741)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3742)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3743)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3744)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3745)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3746)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3747)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3748)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3749)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3750)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3751)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3752)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3753)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3754)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3755)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3756)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3757)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3758)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3759)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3760)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3761)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3762)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3763)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3764)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3765)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3766)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3767)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3768)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3769)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3770)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3771)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3772)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3773)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3774)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3775)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3776)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3777)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3778)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3779)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3780)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3781)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3782)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3783)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3784)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3785)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3786)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3787)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3788)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3789)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3790)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3791)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3792)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3793)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3794)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3795)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3796)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3797)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3798)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3799)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3800)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3801)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3802)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3803)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3804)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3805)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3806)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3807)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3808)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3809)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3810)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3811)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3812)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3813)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3814)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3815)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3816)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3817)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3818)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3819)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3820)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3821)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3822)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3823)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3824)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3825)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3826)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3827)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3828)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3829)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3830)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3831)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3832)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3833)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3834)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3835)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3836)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3837)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3838)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3839)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3840)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3841)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3842)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3843)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3844)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3845)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3846)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3847)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3848)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3849)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3850)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3851)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3852)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3853)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3854)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3855)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3856)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3857)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3858)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3859)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3860)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3861)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3862)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3863)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3864)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3865)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3866)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3867)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3868)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3869)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3870)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3871)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3872)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3873)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3874)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3875)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3876)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3877)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3878)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3879)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3880)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3881)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3882)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3883)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3884)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3885)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3886)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3887)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3888)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3889)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3890)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3891)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3892)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3893)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3894)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3895)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3896)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3897)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3898)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3899)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3900)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3901)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3902)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3903)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3904)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3905)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3906)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3907)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3908)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3909)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3910)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3911)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3912)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3913)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3914)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3915)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3916)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3917)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3918)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3919)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3920)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3921)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3922)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3923)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3924)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3925)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3926)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3927)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3928)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3929)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3930)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3931)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3932)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3933)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3934)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3935)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3936)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3937)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3938)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3939)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(3940)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3941)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3942)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3943)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(3944)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3945)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3946)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3947)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(3948)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3949)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3950)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3951)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(3952)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3953)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3954)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3955)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(3956)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3957)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3958)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3959)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(3960)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3961)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3962)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3963)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(3964)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3965)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3966)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3967)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(3968)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3969)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3970)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3971)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(3972)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3973)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3974)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3975)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(3976)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3977)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3978)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3979)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(3980)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3981)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3982)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3983)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(3984)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3985)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3986)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3987)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(3988)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3989)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3990)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3991)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(3992)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3993)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3994)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3995)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(3996)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3997)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3998)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(3999)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4000)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4001)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4002)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4003)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4004)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4005)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4006)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4007)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4008)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4009)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4010)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4011)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4012)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4013)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4014)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4015)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4016)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4017)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4018)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4019)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4020)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4021)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4022)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4023)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4024)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4025)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4026)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4027)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4028)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4029)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4030)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4031)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4032)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4033)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4034)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4035)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4036)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4037)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4038)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4039)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4040)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4041)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4042)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4043)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4044)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4045)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4046)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4047)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4048)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4049)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4050)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4051)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4052)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4053)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4054)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4055)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4056)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4057)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4058)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4059)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4060)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4061)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4062)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4063)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4064)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4065)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4066)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4067)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4068)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4069)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4070)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4071)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4072)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4073)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4074)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4075)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4076)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4077)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4078)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4079)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4080)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4081)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4082)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4083)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4084)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4085)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4086)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4087)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4088)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4089)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4090)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4091)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4092)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4093)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4094)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4095)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4096)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4097)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4098)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4099)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4100)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4101)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4102)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4103)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4104)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4105)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4106)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4107)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4108)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4109)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4110)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4111)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4112)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4113)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4114)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4115)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4116)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4117)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4118)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4119)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4120)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4121)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4122)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4123)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4124)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4125)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4126)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4127)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4128)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4129)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4130)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4131)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4132)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4133)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4134)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4135)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4136)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4137)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4138)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4139)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4140)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4141)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4142)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4143)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4144)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4145)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4146)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4147)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4148)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4149)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4150)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4151)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4152)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4153)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4154)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4155)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4156)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4157)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4158)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4159)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4160)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4161)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4162)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4163)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4164)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4165)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4166)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4167)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4168)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4169)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4170)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4171)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4172)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4173)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4174)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4175)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4176)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4177)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4178)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4179)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4180)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4181)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4182)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4183)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4184)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4185)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4186)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4187)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4188)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4189)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4190)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4191)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4192)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4193)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4194)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4195)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4196)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4197)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4198)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4199)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4200)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4201)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4202)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4203)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4204)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4205)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4206)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4207)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4208)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4209)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4210)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4211)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4212)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4213)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4214)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4215)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4216)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4217)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4218)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4219)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4220)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4221)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4222)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4223)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4224)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4225)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4226)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4227)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4228)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4229)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4230)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4231)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4232)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4233)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4234)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4235)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4236)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4237)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4238)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4239)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4240)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4241)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4242)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4243)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4244)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4245)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4246)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4247)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4248)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4249)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4250)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4251)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4252)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4253)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4254)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4255)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4256)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4257)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4258)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4259)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4260)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4261)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4262)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4263)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4264)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4265)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4266)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4267)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4268)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4269)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4270)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4271)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4272)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4273)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4274)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4275)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4276)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4277)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4278)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4279)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4280)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4281)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4282)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4283)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4284)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4285)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4286)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4287)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4288)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4289)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4290)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4291)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4292)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4293)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4294)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4295)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4296)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4297)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4298)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4299)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4300)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4301)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4302)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4303)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4304)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4305)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4306)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4307)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4308)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4309)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4310)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4311)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4312)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4313)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4314)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4315)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4316)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4317)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4318)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4319)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4320)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4321)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4322)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4323)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4324)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4325)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4326)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4327)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4328)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4329)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4330)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4331)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4332)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4333)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4334)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4335)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4336)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4337)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4338)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4339)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4340)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4341)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4342)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4343)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4344)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4345)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4346)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4347)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4348)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4349)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4350)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4351)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4352)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4353)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4354)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4355)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4356)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4357)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4358)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4359)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4360)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4361)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4362)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4363)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4364)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4365)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4366)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4367)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4368)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4369)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4370)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4371)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4372)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4373)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4374)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4375)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4376)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4377)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4378)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4379)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4380)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4381)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4382)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4383)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4384)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4385)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4386)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4387)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4388)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4389)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4390)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4391)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4392)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4393)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4394)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4395)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4396)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4397)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4398)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4399)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4400)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4401)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4402)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4403)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4404)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4405)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4406)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4407)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4408)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4409)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4410)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4411)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4412)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4413)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4414)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4415)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4416)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4417)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4418)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4419)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4420)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4421)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4422)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4423)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4424)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4425)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4426)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4427)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4428)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4429)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4430)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4431)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4432)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4433)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4434)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4435)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4436)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4437)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4438)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4439)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4440)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4441)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4442)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4443)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4444)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4445)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4446)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4447)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4448)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4449)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4450)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4451)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4452)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4453)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4454)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4455)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4456)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4457)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4458)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4459)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4460)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4461)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4462)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4463)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4464)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4465)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4466)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4467)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4468)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4469)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4470)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4471)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4472)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4473)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4474)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4475)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4476)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4477)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4478)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4479)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4480)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4481)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4482)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4483)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4484)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4485)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4486)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4487)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4488)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4489)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4490)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4491)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4492)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4493)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4494)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4495)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4496)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4497)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4498)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4499)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4500)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4501)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4502)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4503)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4504)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4505)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4506)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4507)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4508)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4509)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4510)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4511)   <="00000000000000000000000000000000";    --TBD:7
    
	-- xx/xx/xx/xx/xx/xx/xx/xx
    -- xx/xx/xx/ IOUT / IIN / YOUT / YIN / XOUT 
    -- HLT / MEMADDRIN / RAMIN / RAMOUT / INSTOUT / INSTIN / AIN / AOUT 
    -- SUMOUT / SUBTRACT / XIN / OUTREGIN / COUNTEN (PC++) / COUNTOUT (PC) / JUMP(set PC) / FI   
    
    --STAA (8D)
    rom_block(4512)   <="00000000000000000100000000000100";    --STAA:0
    rom_block(4513)   <="00000000000000000100000000000100";    --STAA:0
    rom_block(4514)   <="00000000000000000100000000000100";    --STAA:0
    rom_block(4515)   <="00000000000000000100000000000100";    --STAA:0
    rom_block(4516)   <="00000000000000000001010000001000";    --STAA:1
    rom_block(4517)   <="00000000000000000001010000001000";    --STAA:1
    rom_block(4518)   <="00000000000000000001010000001000";    --STAA:1
    rom_block(4519)   <="00000000000000000001010000001000";    --STAA:1
    rom_block(4520)   <=B"00000000_00000000_01000000_00000100";    --STAA:2
    rom_block(4521)   <=B"00000000_00000000_01000000_00000100";    --STAA:2
    rom_block(4522)   <=B"00000000_00000000_01000000_00000100";    --STAA:2
    rom_block(4523)   <=B"00000000_00000000_01000000_00000100";    --STAA:2
    rom_block(4524)   <=B"00000000_00000000_01010000_00001000";    --STAA:3
    rom_block(4525)   <=B"00000000_00000000_01010000_00001000";    --STAA:3
    rom_block(4526)   <=B"00000000_00000000_01010000_00001000";    --STAA:3
    rom_block(4527)   <=B"00000000_00000000_01010000_00001000";    --STAA:3
    rom_block(4528)   <=B"00000000_00000000_00100001_00000000";    --STAA:4
    rom_block(4529)   <=B"00000000_00000000_00100001_00000000";    --STAA:4
    rom_block(4530)   <=B"00000000_00000000_00100001_00000000";    --STAA:4
    rom_block(4531)   <=B"00000000_00000000_00100001_00000000";    --STAA:4
    rom_block(4532)   <="00000000000000000000000000000000";    --STAA:5
    rom_block(4533)   <="00000000000000000000000000000000";    --STAA:5
    rom_block(4534)   <="00000000000000000000000000000000";    --STAA:5
    rom_block(4535)   <="00000000000000000000000000000000";    --STAA:5
    rom_block(4536)   <="00000000000000000000000000000000";    --STAA:6
    rom_block(4537)   <="00000000000000000000000000000000";    --STAA:6
    rom_block(4538)   <="00000000000000000000000000000000";    --STAA:6
    rom_block(4539)   <="00000000000000000000000000000000";    --STAA:6
    rom_block(4540)   <="00000000000000000000000000000000";    --STAA:7
    rom_block(4541)   <="00000000000000000000000000000000";    --STAA:7
    rom_block(4542)   <="00000000000000000000000000000000";    --STAA:7
    rom_block(4543)   <="00000000000000000000000000000000";    --STAA:7
    
    
    rom_block(4544)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4545)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4546)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4547)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4548)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4549)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4550)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4551)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4552)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4553)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4554)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4555)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4556)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4557)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4558)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4559)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4560)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4561)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4562)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4563)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4564)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4565)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4566)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4567)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4568)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4569)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4570)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4571)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4572)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4573)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4574)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4575)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4576)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4577)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4578)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4579)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4580)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4581)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4582)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4583)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4584)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4585)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4586)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4587)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4588)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4589)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4590)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4591)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4592)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4593)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4594)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4595)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4596)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4597)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4598)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4599)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4600)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4601)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4602)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4603)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4604)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4605)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4606)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4607)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4608)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4609)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4610)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4611)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4612)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4613)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4614)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4615)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4616)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4617)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4618)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4619)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4620)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4621)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4622)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4623)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4624)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4625)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4626)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4627)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4628)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4629)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4630)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4631)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4632)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4633)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4634)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4635)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4636)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4637)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4638)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4639)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4640)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4641)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4642)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4643)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4644)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4645)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4646)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4647)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4648)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4649)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4650)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4651)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4652)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4653)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4654)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4655)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4656)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4657)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4658)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4659)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4660)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4661)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4662)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4663)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4664)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4665)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4666)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4667)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4668)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4669)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4670)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4671)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4672)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4673)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4674)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4675)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4676)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4677)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4678)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4679)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4680)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4681)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4682)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4683)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4684)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4685)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4686)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4687)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4688)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4689)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4690)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4691)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4692)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4693)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4694)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4695)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4696)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4697)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4698)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4699)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4700)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4701)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4702)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4703)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4704)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4705)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4706)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4707)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4708)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4709)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4710)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4711)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4712)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4713)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4714)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4715)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4716)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4717)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4718)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4719)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4720)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4721)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4722)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4723)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4724)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4725)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4726)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4727)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4728)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4729)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4730)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4731)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4732)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4733)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4734)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4735)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4736)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4737)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4738)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4739)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4740)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4741)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4742)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4743)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4744)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4745)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4746)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4747)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4748)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4749)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4750)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4751)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4752)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4753)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4754)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4755)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4756)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4757)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4758)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4759)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4760)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4761)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4762)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4763)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4764)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4765)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4766)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4767)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4768)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4769)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4770)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4771)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4772)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4773)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4774)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4775)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4776)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4777)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4778)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4779)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4780)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4781)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4782)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4783)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4784)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4785)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4786)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4787)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4788)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4789)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4790)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4791)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4792)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4793)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4794)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4795)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4796)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4797)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4798)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4799)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4800)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4801)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4802)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4803)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4804)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4805)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4806)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4807)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4808)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4809)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4810)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4811)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4812)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4813)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4814)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4815)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4816)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4817)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4818)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4819)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4820)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4821)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4822)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4823)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4824)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4825)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4826)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4827)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4828)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4829)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4830)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4831)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4832)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4833)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4834)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4835)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4836)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4837)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4838)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4839)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4840)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4841)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4842)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4843)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4844)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4845)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4846)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4847)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4848)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4849)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4850)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4851)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4852)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4853)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4854)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4855)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4856)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4857)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4858)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4859)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4860)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4861)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4862)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4863)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4864)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4865)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4866)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4867)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4868)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4869)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4870)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4871)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4872)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4873)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4874)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4875)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4876)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4877)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4878)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4879)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4880)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4881)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4882)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4883)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4884)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4885)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4886)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4887)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4888)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4889)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4890)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4891)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4892)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4893)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4894)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4895)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4896)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4897)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4898)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4899)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4900)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4901)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4902)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4903)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4904)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4905)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4906)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4907)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4908)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4909)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4910)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4911)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4912)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4913)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4914)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4915)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4916)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4917)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4918)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4919)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4920)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4921)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4922)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4923)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4924)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4925)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4926)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4927)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4928)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4929)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4930)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4931)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4932)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4933)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4934)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4935)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4936)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4937)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4938)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4939)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(4940)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4941)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4942)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4943)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(4944)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4945)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4946)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4947)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(4948)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4949)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4950)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4951)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(4952)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4953)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4954)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4955)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(4956)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4957)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4958)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4959)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(4960)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4961)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4962)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4963)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(4964)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4965)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4966)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4967)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(4968)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4969)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4970)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4971)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(4972)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4973)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4974)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4975)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(4976)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4977)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4978)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4979)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(4980)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4981)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4982)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4983)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(4984)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4985)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4986)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4987)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(4988)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4989)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4990)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4991)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(4992)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4993)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4994)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4995)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(4996)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4997)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4998)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(4999)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5000)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5001)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5002)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5003)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5004)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5005)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5006)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5007)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5008)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5009)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5010)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5011)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5012)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5013)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5014)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5015)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5016)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5017)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5018)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5019)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5020)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5021)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5022)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5023)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5024)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5025)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5026)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5027)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5028)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5029)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5030)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5031)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5032)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5033)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5034)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5035)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5036)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5037)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5038)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5039)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5040)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5041)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5042)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5043)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5044)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5045)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5046)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5047)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5048)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5049)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5050)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5051)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5052)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5053)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5054)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5055)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5056)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5057)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5058)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5059)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5060)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5061)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5062)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5063)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5064)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5065)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5066)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5067)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5068)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5069)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5070)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5071)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5072)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5073)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5074)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5075)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5076)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5077)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5078)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5079)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5080)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5081)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5082)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5083)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5084)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5085)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5086)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5087)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5088)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5089)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5090)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5091)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5092)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5093)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5094)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5095)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5096)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5097)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5098)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5099)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5100)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5101)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5102)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5103)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5104)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5105)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5106)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5107)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5108)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5109)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5110)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5111)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5112)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5113)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5114)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5115)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5116)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5117)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5118)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5119)   <="00000000000000000000000000000000";    --TBD2:7
    
	-- xx/xx/xx/xx/xx/xx/xx/xx
    -- xx/xx/xx/ IOUT / IIN / YOUT / YIN / XOUT 
    -- HLT / MEMADDRIN / RAMIN / RAMOUT / INSTOUT / INSTIN / AIN / AOUT 
    -- SUMOUT / SUBTRACT / XIN / OUTREGIN / COUNTEN (PC++) / COUNTOUT (PC) / JUMP(set PC) / FI   

    --LDY Immed (A0)
    rom_block(5120)   <="00000000000000000100000000000100";    --LDYI:0             -step 0
    rom_block(5121)   <="00000000000000000100000000000100";    --LDYI:0
    rom_block(5122)   <="00000000000000000100000000000100";    --LDYI:0
    rom_block(5123)   <="00000000000000000100000000000100";    --LDYI:0
    rom_block(5124)   <="00000000000000000001010000001000";    --LDYI:1             -step 1
    rom_block(5125)   <="00000000000000000001010000001000";    --LDYI:1
    rom_block(5126)   <="00000000000000000001010000001000";    --LDYI:1
    rom_block(5127)   <="00000000000000000001010000001000";    --LDYI:1
    rom_block(5128)   <="00000000000000000100000000000100";    --LDYI:2             -step 2                 
    rom_block(5129)   <="00000000000000000100000000000100";    --LDYI:2
    rom_block(5130)   <="00000000000000000100000000000100";    --LDYI:2
    rom_block(5131)   <="00000000000000000100000000000100";    --LDYI:2
    rom_block(5132)   <="00000000000000100001000000001000";    --LDYI:3
    rom_block(5133)   <=B"0000000000000010_0001000000001000";    --LDYI:3
    rom_block(5134)   <=B"0000000000000010_0001000000001000";    --LDYI:3
    rom_block(5135)   <=B"0000000000000010_0001000000001000";    --LDYI:3
    rom_block(5136)   <=B"0000000000000000_0000000000000100";    --LDYI:4
    rom_block(5137)   <="00000000000000000000000000000100";    --LDYI:4
    rom_block(5138)   <="00000000000000000000000000000100";    --LDYI:4
    rom_block(5139)   <="00000000000000000000000000000100";    --LDYI:4
    rom_block(5140)   <="00000000000000000000000000000000";    --LDYI:5
    rom_block(5141)   <="00000000000000000000000000000000";    --LDYI:5
    rom_block(5142)   <="00000000000000000000000000000000";    --LDYI:5
    rom_block(5143)   <="00000000000000000000000000000000";    --LDYI:5
    rom_block(5144)   <="00000000000000000000000000000000";    --LDYI:6
    rom_block(5145)   <="00000000000000000000000000000000";    --LDYI:6
    rom_block(5146)   <="00000000000000000000000000000000";    --LDYI:6
    rom_block(5147)   <="00000000000000000000000000000000";    --LDYI:6
    rom_block(5148)   <="00000000000000000000000000000000";    --LDYI:7
    rom_block(5149)   <="00000000000000000000000000000000";    --LDYI:7
    rom_block(5150)   <="00000000000000000000000000000000";    --LDYI:7
    rom_block(5151)   <="00000000000000000000000000000000";    --LDYI:7
    
    rom_block(5152)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5153)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5154)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5155)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5156)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5157)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5158)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5159)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5160)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5161)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5162)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5163)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5164)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5165)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5166)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5167)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5168)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5169)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5170)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5171)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5172)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5173)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5174)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5175)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5176)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5177)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5178)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5179)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5180)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5181)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5182)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5183)   <="00000000000000000000000000000000";    --TBD2:7
    
    -- IOUT / IIN / YOUT / YIN / XOUT / HLT / MEMADDRIN / RAMIN / RAMOUT / INSTOUT / INSTIN / AIN / AOUT / SUMOUT / SUBTRACT / XIN / OUTREGIN / COUNTEN (PC++) / COUNTOUT (PC) / JUMP(set PC) / FI
    --LDX Immed (A2)
    rom_block(5184)   <="00000000000000000100000000000100";    --LDXI:0
    rom_block(5185)   <="00000000000000000100000000000100";    --LDXI:0
    rom_block(5186)   <="00000000000000000100000000000100";    --LDXI:0
    rom_block(5187)   <="00000000000000000100000000000100";    --LDXI:0
    rom_block(5188)   <="00000000000000000001010000001000";    --LDXI:1
    rom_block(5189)   <="00000000000000000001010000001000";    --LDXI:1
    rom_block(5190)   <="00000000000000000001010000001000";    --LDXI:1
    rom_block(5191)   <="00000000000000000001010000001000";    --LDXI:1
    rom_block(5192)   <="00000000000000000100000000000100";    --LDXI:2
    rom_block(5193)   <="00000000000000000100000000000100";    --LDXI:2
    rom_block(5194)   <="00000000000000000100000000000100";    --LDXI:2
    rom_block(5195)   <="00000000000000000100000000000100";    --LDXI:2
    rom_block(5196)   <="00000000000000000001000000101000";    --LDXI:3
    rom_block(5197)   <="00000000000000000001000000101000";    --LDXI:3
    rom_block(5198)   <="00000000000000000001000000101000";    --LDXI:3
    rom_block(5199)   <="00000000000000000001000000101000";    --LDXI:3
    rom_block(5200)   <="00000000000000000000000000000100";    --LDXI:4
    rom_block(5201)   <="00000000000000000000000000000100";    --LDXI:4
    rom_block(5202)   <="00000000000000000000000000000100";    --LDXI:4
    rom_block(5203)   <="00000000000000000000000000000100";    --LDXI:4
    rom_block(5204)   <="00000000000000000000000000000000";    --LDXI:5
    rom_block(5205)   <="00000000000000000000000000000000";    --LDXI:5
    rom_block(5206)   <="00000000000000000000000000000000";    --LDXI:5
    rom_block(5207)   <="00000000000000000000000000000000";    --LDXI:5
    rom_block(5208)   <="00000000000000000000000000000000";    --LDXI:6
    rom_block(5209)   <="00000000000000000000000000000000";    --LDXI:6
    rom_block(5210)   <="00000000000000000000000000000000";    --LDXI:6
    rom_block(5211)   <="00000000000000000000000000000000";    --LDXI:6
    rom_block(5212)   <="00000000000000000000000000000000";    --LDXI:7
    rom_block(5213)   <="00000000000000000000000000000000";    --LDXI:7
    rom_block(5214)   <="00000000000000000000000000000000";    --LDXI:7
    rom_block(5215)   <="00000000000000000000000000000000";    --LDXI:7
    
    rom_block(5216)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5217)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5218)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5219)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5220)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5221)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5222)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5223)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5224)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5225)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5226)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5227)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5228)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5229)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5230)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5231)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5232)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5233)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5234)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5235)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5236)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5237)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5238)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5239)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5240)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5241)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5242)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5243)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5244)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5245)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5246)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5247)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5248)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5249)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5250)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5251)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5252)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5253)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5254)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5255)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5256)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5257)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5258)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5259)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5260)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5261)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5262)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5263)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5264)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5265)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5266)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5267)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5268)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5269)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5270)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5271)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5272)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5273)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5274)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5275)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5276)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5277)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5278)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5279)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5280)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5281)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5282)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5283)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5284)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5285)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5286)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5287)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5288)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5289)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5290)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5291)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5292)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5293)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5294)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5295)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5296)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5297)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5298)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5299)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5300)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5301)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5302)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5303)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5304)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5305)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5306)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5307)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5308)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5309)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5310)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5311)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5312)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5313)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5314)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5315)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5316)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5317)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5318)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5319)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5320)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5321)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5322)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5323)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5324)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5325)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5326)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5327)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5328)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5329)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5330)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5331)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5332)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5333)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5334)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5335)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5336)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5337)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5338)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5339)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5340)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5341)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5342)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5343)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5344)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5345)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5346)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5347)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5348)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5349)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5350)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5351)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5352)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5353)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5354)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5355)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5356)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5357)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5358)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5359)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5360)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5361)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5362)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5363)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5364)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5365)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5366)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5367)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5368)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5369)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5370)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5371)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5372)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5373)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5374)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5375)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5376)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5377)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5378)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5379)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5380)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5381)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5382)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5383)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5384)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5385)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5386)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5387)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5388)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5389)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5390)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5391)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5392)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5393)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5394)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5395)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5396)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5397)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5398)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5399)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5400)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5401)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5402)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5403)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5404)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5405)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5406)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5407)   <="00000000000000000000000000000000";    --TBD:7

	-- xx/xx/xx/xx/xx/xx/xx/xx
    -- xx/xx/xx/ IOUT / IIN / YOUT / YIN / XOUT 
    -- HLT / MEMADDRIN / RAMIN / RAMOUT / INSTOUT / INSTIN / AIN / AOUT 
    -- SUMOUT / SUBTRACT / XIN / OUTREGIN / COUNTEN (PC++) / COUNTOUT (PC) / JUMP(set PC) / FI   

--    --LDA Immediate (A9)
    rom_block(5408)   <="00000000000000000100000000000100";    --LDAI:0             -step 0
    rom_block(5409)   <="00000000000000000100000000000100";    --LDAI:0
    rom_block(5410)   <="00000000000000000100000000000100";    --LDAI:0
    rom_block(5411)   <="00000000000000000100000000000100";    --LDAI:0
    rom_block(5412)   <="00000000000000000001010000001000";    --LDAI:1             -step 1
    rom_block(5413)   <="00000000000000000001010000001000";    --LDAI:1
    rom_block(5414)   <="00000000000000000001010000001000";    --LDAI:1
    rom_block(5415)   <="00000000000000000001010000001000";    --LDAI:1
    rom_block(5416)   <=B"00000000_00000000_01000000_00000100";    --LDAI:2             -step 2                 
    rom_block(5417)   <=B"00000000_00000000_01000000_00000100";    --LDAI:2
    rom_block(5418)   <=B"00000000_00000000_01000000_00000100";    --LDAI:2
    rom_block(5419)   <=B"00000000_00000000_01000000_00000100";    --LDAI:2
    rom_block(5420)   <=B"00000000_00000000_00010010_00001000";    --LDAI:3
    rom_block(5421)   <=B"00000000_00000000_00010010_00001000";    --LDAI:3
    rom_block(5422)   <=B"00000000_00000000_00010010_00001000";    --LDAI:3
    rom_block(5423)   <=B"00000000_00000000_00010010_00001000";    --LDAI:3
    rom_block(5424)   <="00000000000000000000000000000100";    --LDAI:4
    rom_block(5425)   <="00000000000000000000000000000100";    --LDAI:4
    rom_block(5426)   <="00000000000000000000000000000100";    --LDAI:4
    rom_block(5427)   <="00000000000000000000000000000100";    --LDAI:4
    rom_block(5428)   <="00000000000000000000000000000000";    --LDAI:5
    rom_block(5429)   <="00000000000000000000000000000000";    --LDAI:5
    rom_block(5430)   <="00000000000000000000000000000000";    --LDAI:5
    rom_block(5431)   <="00000000000000000000000000000000";    --LDAI:5
    rom_block(5432)   <="00000000000000000000000000000000";    --LDAI:6
    rom_block(5433)   <="00000000000000000000000000000000";    --LDAI:6
    rom_block(5434)   <="00000000000000000000000000000000";    --LDAI:6
    rom_block(5435)   <="00000000000000000000000000000000";    --LDAI:6
    rom_block(5436)   <="00000000000000000000000000000000";    --LDAI:7
    rom_block(5437)   <="00000000000000000000000000000000";    --LDAI:7
    rom_block(5438)   <="00000000000000000000000000000000";    --LDAI:7
    rom_block(5439)   <="00000000000000000000000000000000";    --LDAI:7
    
    rom_block(5440)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5441)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5442)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5443)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5444)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5445)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5446)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5447)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5448)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5449)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5450)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5451)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5452)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5453)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5454)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5455)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5456)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5457)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5458)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5459)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5460)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5461)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5462)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5463)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5464)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5465)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5466)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5467)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5468)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5469)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5470)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5471)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5472)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5473)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5474)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5475)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5476)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5477)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5478)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5479)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5480)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5481)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5482)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5483)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5484)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5485)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5486)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5487)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5488)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5489)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5490)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5491)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5492)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5493)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5494)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5495)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5496)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5497)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5498)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5499)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5500)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5501)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5502)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5503)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5504)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5505)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5506)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5507)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5508)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5509)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5510)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5511)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5512)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5513)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5514)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5515)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5516)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5517)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5518)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5519)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5520)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5521)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5522)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5523)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5524)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5525)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5526)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5527)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5528)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5529)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5530)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5531)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5532)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5533)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5534)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5535)   <="00000000000000000000000000000000";    --TBD:7
    
    --LDAA (AD)
    rom_block(5536)   <="00000000000000000100000000000100";    --LDAA:0
    rom_block(5537)   <="00000000000000000100000000000100";    --LDAA:0
    rom_block(5538)   <="00000000000000000100000000000100";    --LDAA:0
    rom_block(5539)   <="00000000000000000100000000000100";    --LDAA:0
    rom_block(5540)   <="00000000000000000001010000001000";    --LDAA:1
    rom_block(5541)   <="00000000000000000001010000001000";    --LDAA:1
    rom_block(5542)   <="00000000000000000001010000001000";    --LDAA:1
    rom_block(5543)   <="00000000000000000001010000001000";    --LDAA:1
    rom_block(5544)   <="00000000000000000100000000000100";    --LDAA:2
    rom_block(5545)   <="00000000000000000100000000000100";    --LDAA:2
    rom_block(5546)   <="00000000000000000100000000000100";    --LDAA:2
    rom_block(5547)   <="00000000000000000100000000000100";    --LDAA:2
    rom_block(5548)   <="00000000000000000101000000001000";    --LDAA:3
    rom_block(5549)   <="00000000000000000101000000001000";    --LDAA:3
    rom_block(5550)   <="00000000000000000101000000001000";    --LDAA:3
    rom_block(5551)   <="00000000000000000101000000001000";    --LDAA:3
    rom_block(5552)   <="00000000000000000001001000000000";    --LDAA:4
    rom_block(5553)   <="00000000000000000001001000000000";    --LDAA:4
    rom_block(5554)   <="00000000000000000001001000000000";    --LDAA:4
    rom_block(5555)   <="00000000000000000001001000000000";    --LDAA:4
    rom_block(5556)   <="00000000000000000000000000000000";    --LDAA:5
    rom_block(5557)   <="00000000000000000000000000000000";    --LDAA:5
    rom_block(5558)   <="00000000000000000000000000000000";    --LDAA:5
    rom_block(5559)   <="00000000000000000000000000000000";    --LDAA:5
    rom_block(5560)   <="00000000000000000000000000000000";    --LDAA:6
    rom_block(5561)   <="00000000000000000000000000000000";    --LDAA:6
    rom_block(5562)   <="00000000000000000000000000000000";    --LDAA:6
    rom_block(5563)   <="00000000000000000000000000000000";    --LDAA:6
    rom_block(5564)   <="00000000000000000000000000000000";    --LDAA:7
    rom_block(5565)   <="00000000000000000000000000000000";    --LDAA:7
    rom_block(5566)   <="00000000000000000000000000000000";    --LDAA:7
    rom_block(5567)   <="00000000000000000000000000000000";    --LDAA:7
    
    rom_block(5568)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5569)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5570)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5571)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5572)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5573)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5574)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5575)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5576)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5577)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5578)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5579)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5580)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5581)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5582)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5583)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5584)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5585)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5586)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5587)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5588)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5589)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5590)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5591)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5592)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5593)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5594)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5595)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5596)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5597)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5598)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5599)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5600)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5601)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5602)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5603)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5604)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5605)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5606)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5607)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5608)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5609)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5610)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5611)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5612)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5613)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5614)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5615)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5616)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5617)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5618)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5619)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5620)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5621)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5622)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5623)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5624)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5625)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5626)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5627)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5628)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5629)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5630)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5631)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5632)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5633)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5634)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5635)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5636)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5637)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5638)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5639)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5640)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5641)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5642)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5643)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5644)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5645)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5646)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5647)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5648)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5649)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5650)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5651)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5652)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5653)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5654)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5655)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5656)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5657)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5658)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5659)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5660)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5661)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5662)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5663)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5664)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5665)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5666)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5667)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5668)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5669)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5670)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5671)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5672)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5673)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5674)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5675)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5676)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5677)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5678)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5679)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5680)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5681)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5682)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5683)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5684)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5685)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5686)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5687)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5688)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5689)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5690)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5691)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5692)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5693)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5694)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5695)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5696)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5697)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5698)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5699)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5700)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5701)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5702)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5703)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5704)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5705)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5706)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5707)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5708)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5709)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5710)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5711)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5712)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5713)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5714)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5715)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5716)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5717)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5718)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5719)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5720)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5721)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5722)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5723)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5724)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5725)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5726)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5727)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5728)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5729)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5730)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5731)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5732)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5733)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5734)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5735)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5736)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5737)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5738)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5739)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5740)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5741)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5742)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5743)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5744)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5745)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5746)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5747)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5748)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5749)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5750)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5751)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5752)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5753)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5754)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5755)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5756)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5757)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5758)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5759)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5760)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5761)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5762)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5763)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5764)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5765)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5766)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5767)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5768)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5769)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5770)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5771)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5772)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5773)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5774)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5775)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5776)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5777)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5778)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5779)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5780)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5781)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5782)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5783)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5784)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5785)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5786)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5787)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5788)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5789)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5790)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5791)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5792)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5793)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5794)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5795)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5796)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5797)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5798)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5799)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5800)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5801)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5802)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5803)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5804)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5805)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5806)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5807)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5808)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5809)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5810)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5811)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5812)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5813)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5814)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5815)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5816)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5817)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5818)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5819)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5820)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5821)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5822)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5823)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5824)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5825)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5826)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5827)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5828)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5829)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5830)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5831)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5832)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5833)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5834)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5835)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5836)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5837)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5838)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5839)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5840)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5841)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5842)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5843)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5844)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5845)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5846)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5847)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5848)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5849)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5850)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5851)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5852)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5853)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5854)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5855)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5856)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5857)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5858)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5859)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5860)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5861)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5862)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5863)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5864)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5865)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5866)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5867)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5868)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5869)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5870)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5871)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5872)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5873)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5874)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5875)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5876)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5877)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5878)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5879)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5880)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5881)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5882)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5883)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5884)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5885)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5886)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5887)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5888)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5889)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5890)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5891)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5892)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5893)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5894)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5895)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5896)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5897)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5898)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5899)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5900)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5901)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5902)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5903)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5904)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5905)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5906)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5907)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5908)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5909)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5910)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5911)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5912)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5913)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5914)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5915)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5916)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5917)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5918)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5919)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5920)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5921)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5922)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5923)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5924)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5925)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5926)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5927)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5928)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5929)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5930)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5931)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5932)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5933)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5934)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5935)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5936)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5937)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5938)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5939)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(5940)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5941)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5942)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5943)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(5944)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5945)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5946)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5947)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(5948)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5949)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5950)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5951)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(5952)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5953)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5954)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5955)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(5956)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5957)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5958)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5959)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(5960)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5961)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5962)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5963)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(5964)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5965)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5966)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5967)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(5968)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5969)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5970)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5971)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(5972)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5973)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5974)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5975)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(5976)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5977)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5978)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5979)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(5980)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5981)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5982)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5983)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(5984)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5985)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5986)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5987)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(5988)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5989)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5990)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5991)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(5992)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5993)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5994)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5995)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(5996)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5997)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5998)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(5999)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6000)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6001)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6002)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6003)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6004)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6005)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6006)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6007)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6008)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6009)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6010)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6011)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6012)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6013)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6014)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6015)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6016)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6017)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6018)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6019)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6020)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6021)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6022)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6023)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6024)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6025)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6026)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6027)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6028)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6029)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6030)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6031)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6032)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6033)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6034)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6035)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6036)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6037)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6038)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6039)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6040)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6041)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6042)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6043)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6044)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6045)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6046)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6047)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6048)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6049)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6050)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6051)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6052)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6053)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6054)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6055)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6056)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6057)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6058)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6059)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6060)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6061)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6062)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6063)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6064)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6065)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6066)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6067)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6068)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6069)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6070)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6071)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6072)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6073)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6074)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6075)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6076)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6077)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6078)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6079)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6080)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6081)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6082)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6083)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6084)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6085)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6086)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6087)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6088)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6089)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6090)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6091)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6092)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6093)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6094)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6095)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6096)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6097)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6098)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6099)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6100)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6101)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6102)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6103)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6104)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6105)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6106)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6107)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6108)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6109)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6110)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6111)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6112)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6113)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6114)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6115)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6116)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6117)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6118)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6119)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6120)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6121)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6122)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6123)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6124)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6125)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6126)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6127)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6128)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6129)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6130)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6131)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6132)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6133)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6134)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6135)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6136)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6137)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6138)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6139)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6140)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6141)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6142)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6143)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6144)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6145)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6146)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6147)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6148)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6149)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6150)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6151)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6152)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6153)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6154)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6155)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6156)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6157)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6158)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6159)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6160)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6161)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6162)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6163)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6164)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6165)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6166)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6167)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6168)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6169)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6170)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6171)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6172)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6173)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6174)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6175)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6176)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6177)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6178)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6179)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6180)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6181)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6182)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6183)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6184)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6185)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6186)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6187)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6188)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6189)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6190)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6191)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6192)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6193)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6194)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6195)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6196)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6197)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6198)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6199)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6200)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6201)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6202)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6203)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6204)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6205)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6206)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6207)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6208)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6209)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6210)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6211)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6212)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6213)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6214)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6215)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6216)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6217)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6218)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6219)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6220)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6221)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6222)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6223)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6224)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6225)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6226)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6227)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6228)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6229)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6230)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6231)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6232)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6233)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6234)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6235)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6236)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6237)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6238)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6239)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6240)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6241)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6242)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6243)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6244)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6245)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6246)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6247)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6248)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6249)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6250)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6251)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6252)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6253)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6254)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6255)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6256)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6257)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6258)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6259)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6260)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6261)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6262)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6263)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6264)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6265)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6266)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6267)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6268)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6269)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6270)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6271)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6272)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6273)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6274)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6275)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6276)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6277)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6278)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6279)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6280)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6281)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6282)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6283)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6284)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6285)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6286)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6287)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6288)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6289)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6290)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6291)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6292)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6293)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6294)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6295)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6296)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6297)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6298)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6299)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6300)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6301)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6302)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6303)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6304)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6305)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6306)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6307)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6308)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6309)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6310)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6311)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6312)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6313)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6314)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6315)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6316)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6317)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6318)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6319)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6320)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6321)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6322)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6323)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6324)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6325)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6326)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6327)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6328)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6329)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6330)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6331)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6332)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6333)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6334)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6335)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6336)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6337)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6338)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6339)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6340)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6341)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6342)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6343)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6344)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6345)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6346)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6347)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6348)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6349)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6350)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6351)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6352)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6353)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6354)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6355)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6356)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6357)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6358)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6359)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6360)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6361)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6362)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6363)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6364)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6365)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6366)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6367)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6368)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6369)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6370)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6371)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6372)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6373)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6374)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6375)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6376)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6377)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6378)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6379)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6380)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6381)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6382)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6383)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6384)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6385)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6386)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6387)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6388)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6389)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6390)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6391)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6392)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6393)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6394)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6395)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6396)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6397)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6398)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6399)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6400)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6401)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6402)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6403)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6404)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6405)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6406)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6407)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6408)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6409)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6410)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6411)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6412)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6413)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6414)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6415)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6416)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6417)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6418)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6419)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6420)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6421)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6422)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6423)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6424)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6425)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6426)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6427)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6428)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6429)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6430)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6431)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6432)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6433)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6434)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6435)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6436)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6437)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6438)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6439)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6440)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6441)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6442)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6443)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6444)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6445)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6446)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6447)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6448)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6449)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6450)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6451)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6452)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6453)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6454)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6455)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6456)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6457)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6458)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6459)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6460)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6461)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6462)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6463)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6464)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6465)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6466)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6467)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6468)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6469)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6470)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6471)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6472)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6473)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6474)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6475)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6476)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6477)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6478)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6479)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6480)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6481)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6482)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6483)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6484)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6485)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6486)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6487)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6488)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6489)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6490)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6491)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6492)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6493)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6494)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6495)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6496)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6497)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6498)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6499)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6500)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6501)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6502)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6503)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6504)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6505)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6506)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6507)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6508)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6509)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6510)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6511)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6512)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6513)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6514)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6515)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6516)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6517)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6518)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6519)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6520)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6521)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6522)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6523)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6524)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6525)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6526)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6527)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6528)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6529)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6530)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6531)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6532)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6533)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6534)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6535)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6536)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6537)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6538)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6539)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6540)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6541)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6542)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6543)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6544)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6545)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6546)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6547)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6548)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6549)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6550)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6551)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6552)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6553)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6554)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6555)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6556)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6557)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6558)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6559)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6560)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6561)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6562)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6563)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6564)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6565)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6566)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6567)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6568)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6569)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6570)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6571)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6572)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6573)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6574)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6575)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6576)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6577)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6578)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6579)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6580)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6581)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6582)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6583)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6584)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6585)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6586)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6587)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6588)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6589)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6590)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6591)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6592)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6593)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6594)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6595)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6596)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6597)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6598)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6599)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6600)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6601)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6602)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6603)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6604)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6605)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6606)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6607)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6608)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6609)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6610)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6611)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6612)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6613)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6614)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6615)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6616)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6617)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6618)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6619)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6620)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6621)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6622)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6623)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6624)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6625)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6626)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6627)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6628)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6629)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6630)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6631)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6632)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6633)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6634)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6635)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6636)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6637)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6638)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6639)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6640)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6641)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6642)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6643)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6644)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6645)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6646)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6647)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6648)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6649)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6650)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6651)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6652)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6653)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6654)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6655)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6656)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6657)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6658)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6659)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6660)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6661)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6662)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6663)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6664)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6665)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6666)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6667)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6668)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6669)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6670)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6671)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6672)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6673)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6674)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6675)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6676)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6677)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6678)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6679)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6680)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6681)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6682)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6683)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6684)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6685)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6686)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6687)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6688)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6689)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6690)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6691)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6692)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6693)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6694)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6695)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6696)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6697)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6698)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6699)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6700)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6701)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6702)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6703)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6704)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6705)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6706)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6707)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6708)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6709)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6710)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6711)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6712)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6713)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6714)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6715)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6716)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6717)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6718)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6719)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6720)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6721)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6722)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6723)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6724)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6725)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6726)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6727)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6728)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6729)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6730)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6731)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6732)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6733)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6734)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6735)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6736)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6737)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6738)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6739)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6740)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6741)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6742)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6743)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6744)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6745)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6746)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6747)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6748)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6749)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6750)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6751)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6752)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6753)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6754)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6755)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6756)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6757)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6758)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6759)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6760)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6761)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6762)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6763)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6764)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6765)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6766)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6767)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6768)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6769)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6770)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6771)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6772)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6773)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6774)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6775)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6776)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6777)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6778)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6779)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6780)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6781)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6782)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6783)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6784)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6785)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6786)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6787)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6788)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6789)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6790)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6791)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6792)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6793)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6794)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6795)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6796)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6797)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6798)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6799)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6800)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6801)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6802)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6803)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6804)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6805)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6806)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6807)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6808)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6809)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6810)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6811)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6812)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6813)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6814)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6815)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6816)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6817)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6818)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6819)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6820)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6821)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6822)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6823)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6824)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6825)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6826)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6827)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6828)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6829)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6830)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6831)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6832)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6833)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6834)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6835)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6836)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6837)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6838)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6839)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6840)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6841)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6842)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6843)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6844)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6845)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6846)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6847)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6848)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6849)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6850)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6851)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6852)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6853)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6854)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6855)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6856)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6857)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6858)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6859)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6860)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6861)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6862)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6863)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6864)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6865)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6866)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6867)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6868)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6869)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6870)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6871)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6872)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6873)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6874)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6875)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6876)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6877)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6878)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6879)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6880)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6881)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6882)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6883)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6884)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6885)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6886)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6887)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6888)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6889)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6890)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6891)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6892)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6893)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6894)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6895)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6896)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6897)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6898)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6899)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6900)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6901)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6902)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6903)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6904)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6905)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6906)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6907)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6908)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6909)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6910)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6911)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6912)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6913)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6914)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6915)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6916)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6917)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6918)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6919)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6920)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6921)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6922)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6923)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6924)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6925)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6926)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6927)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6928)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6929)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6930)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6931)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6932)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6933)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6934)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6935)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6936)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6937)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6938)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6939)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(6940)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6941)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6942)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6943)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(6944)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6945)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6946)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6947)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(6948)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6949)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6950)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6951)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(6952)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6953)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6954)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6955)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(6956)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6957)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6958)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6959)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(6960)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6961)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6962)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6963)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(6964)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6965)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6966)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6967)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(6968)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6969)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6970)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6971)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(6972)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6973)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6974)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6975)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(6976)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6977)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6978)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6979)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(6980)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6981)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6982)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6983)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(6984)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6985)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6986)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6987)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(6988)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6989)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6990)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6991)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(6992)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6993)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6994)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6995)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(6996)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6997)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6998)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(6999)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7000)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7001)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7002)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7003)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7004)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7005)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7006)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7007)   <="00000000000000000000000000000000";    --TBD:7
    
    --STP (HALT)
    rom_block(7008)   <="00000000000000000100000000000100";    --STP:0
    rom_block(7009)   <="00000000000000000100000000000100";    --STP:0
    rom_block(7010)   <="00000000000000000100000000000100";    --STP:0
    rom_block(7011)   <="00000000000000000100000000000100";    --STP:0
    rom_block(7012)   <="00000000000000000001010000001000";    --STP:1
    rom_block(7013)   <="00000000000000000001010000001000";    --STP:1
    rom_block(7014)   <="00000000000000000001010000001000";    --STP:1
    rom_block(7015)   <="00000000000000000001010000001000";    --STP:1
    rom_block(7016)   <="00000000000000001000000000000000";    --STP:2
    rom_block(7017)   <="00000000000000001000000000000000";    --STP:2
    rom_block(7018)   <="00000000000000001000000000000000";    --STP:2
    rom_block(7019)   <="00000000000000001000000000000000";    --STP:2
    rom_block(7020)   <="00000000000000000000000000000000";    --STP:3
    rom_block(7021)   <="00000000000000000000000000000000";    --STP:3
    rom_block(7022)   <="00000000000000000000000000000000";    --STP:3
    rom_block(7023)   <="00000000000000000000000000000000";    --STP:3
    rom_block(7024)   <="00000000000000000000000000000000";    --STP:4
    rom_block(7025)   <="00000000000000000000000000000000";    --STP:4
    rom_block(7026)   <="00000000000000000000000000000000";    --STP:4
    rom_block(7027)   <="00000000000000000000000000000000";    --STP:4
    rom_block(7028)   <="00000000000000000000000000000000";    --STP:5
    rom_block(7029)   <="00000000000000000000000000000000";    --STP:5
    rom_block(7030)   <="00000000000000000000000000000000";    --STP:5
    rom_block(7031)   <="00000000000000000000000000000000";    --STP:5
    rom_block(7032)   <="00000000000000000000000000000000";    --STP:6
    rom_block(7033)   <="00000000000000000000000000000000";    --STP:6
    rom_block(7034)   <="00000000000000000000000000000000";    --STP:6
    rom_block(7035)   <="00000000000000000000000000000000";    --STP:6
    rom_block(7036)   <="00000000000000000000000000000000";    --STP:7
    rom_block(7037)   <="00000000000000000000000000000000";    --STP:7
    rom_block(7038)   <="00000000000000000000000000000000";    --STP:7
    rom_block(7039)   <="00000000000000000000000000000000";    --STP:7
    rom_block(7040)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7041)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7042)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7043)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7044)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7045)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7046)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7047)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7048)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7049)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7050)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7051)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7052)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7053)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7054)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7055)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7056)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7057)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7058)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7059)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7060)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7061)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7062)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7063)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7064)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7065)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7066)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7067)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7068)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7069)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7070)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7071)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7072)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7073)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7074)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7075)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7076)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7077)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7078)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7079)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7080)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7081)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7082)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7083)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7084)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7085)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7086)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7087)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7088)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7089)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7090)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7091)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7092)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7093)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7094)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7095)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7096)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7097)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7098)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7099)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7100)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7101)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7102)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7103)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7104)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7105)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7106)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7107)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7108)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7109)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7110)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7111)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7112)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7113)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7114)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7115)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7116)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7117)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7118)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7119)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7120)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7121)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7122)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7123)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7124)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7125)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7126)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7127)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7128)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7129)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7130)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7131)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7132)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7133)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7134)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7135)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7136)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7137)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7138)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7139)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7140)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7141)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7142)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7143)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7144)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7145)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7146)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7147)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7148)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7149)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7150)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7151)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7152)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7153)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7154)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7155)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7156)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7157)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7158)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7159)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7160)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7161)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7162)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7163)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7164)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7165)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7166)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7167)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7168)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7169)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7170)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7171)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7172)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7173)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7174)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7175)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7176)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7177)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7178)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7179)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7180)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7181)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7182)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7183)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7184)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7185)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7186)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7187)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7188)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7189)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7190)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7191)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7192)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7193)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7194)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7195)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7196)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7197)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7198)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7199)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7200)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7201)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7202)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7203)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7204)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7205)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7206)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7207)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7208)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7209)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7210)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7211)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7212)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7213)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7214)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7215)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7216)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7217)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7218)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7219)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7220)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7221)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7222)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7223)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7224)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7225)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7226)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7227)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7228)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7229)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7230)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7231)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7232)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7233)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7234)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7235)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7236)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7237)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7238)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7239)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7240)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7241)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7242)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7243)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7244)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7245)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7246)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7247)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7248)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7249)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7250)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7251)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7252)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7253)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7254)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7255)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7256)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7257)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7258)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7259)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7260)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7261)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7262)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7263)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7264)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7265)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7266)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7267)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7268)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7269)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7270)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7271)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7272)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7273)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7274)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7275)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7276)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7277)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7278)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7279)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7280)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7281)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7282)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7283)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7284)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7285)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7286)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7287)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7288)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7289)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7290)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7291)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7292)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7293)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7294)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7295)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7296)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7297)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7298)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7299)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7300)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7301)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7302)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7303)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7304)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7305)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7306)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7307)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7308)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7309)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7310)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7311)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7312)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7313)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7314)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7315)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7316)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7317)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7318)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7319)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7320)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7321)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7322)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7323)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7324)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7325)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7326)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7327)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7328)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7329)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7330)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7331)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7332)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7333)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7334)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7335)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7336)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7337)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7338)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7339)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7340)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7341)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7342)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7343)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7344)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7345)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7346)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7347)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7348)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7349)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7350)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7351)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7352)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7353)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7354)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7355)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7356)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7357)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7358)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7359)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7360)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7361)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7362)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7363)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7364)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7365)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7366)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7367)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7368)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7369)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7370)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7371)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7372)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7373)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7374)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7375)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7376)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7377)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7378)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7379)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7380)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7381)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7382)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7383)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7384)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7385)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7386)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7387)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7388)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7389)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7390)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7391)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7392)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7393)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7394)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7395)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7396)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7397)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7398)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7399)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7400)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7401)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7402)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7403)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7404)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7405)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7406)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7407)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7408)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7409)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7410)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7411)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7412)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7413)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7414)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7415)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7416)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7417)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7418)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7419)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7420)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7421)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7422)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7423)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7424)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7425)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7426)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7427)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7428)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7429)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7430)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7431)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7432)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7433)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7434)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7435)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7436)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7437)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7438)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7439)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7440)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7441)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7442)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7443)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7444)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7445)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7446)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7447)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7448)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7449)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7450)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7451)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7452)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7453)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7454)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7455)   <="00000000000000000000000000000000";    --TBD:7
    
    -- xx/xx/xx/xx/xx/xx/xx/xx
    -- xx/xx/xx/ IOUT / IIN / YOUT / YIN / XOUT 
    -- HLT / MEMADDRIN / RAMIN / RAMOUT / INSTOUT / INSTIN / AIN / AOUT 
    -- SUMOUT / SUBTRACT / XIN / OUTREGIN / COUNTEN (PC++) / COUNTOUT (PC) / JUMP(set PC) / FI   
    
    --SBC Immed (E9)
    rom_block(7456)   <="00000000000000000100000000000100";    --SBCI:0
    rom_block(7457)   <="00000000000000000100000000000100";    --SBCI:0
    rom_block(7458)   <="00000000000000000100000000000100";    --SBCI:0
    rom_block(7459)   <="00000000000000000100000000000100";    --SBCI:0
    rom_block(7460)   <="00000000000000000001010000001000";    --SBCI:1
    rom_block(7461)   <="00000000000000000001010000001000";    --SBCI:1
    rom_block(7462)   <="00000000000000000001010000001000";    --SBCI:1
    rom_block(7463)   <="00000000000000000001010000001000";    --SBCI:1
    rom_block(7464)   <=B"0000000000000000_0100000000000100";    --SBCI:2
    rom_block(7465)   <=B"0000000000000000_0100000000000100";    --SBCI:2
    rom_block(7466)   <=B"0000000000000000_0100000000000100";    --SBCI:2
    rom_block(7467)   <=B"0000000000000000_0100000000000100";    --SBCI:2
    rom_block(7468)   <=B"0000000000001000_0001000000001000";    --SBCI:3
    rom_block(7469)   <=B"0000000000001000_0001000000001000";    --SBCI:3
    rom_block(7470)   <=B"0000000000001000_0001000000001000";    --SBCI:3
    rom_block(7471)   <=B"0000000000001000_0001000000001000";    --SBCI:3
    rom_block(7472)   <=B"0000000000000000_00000010_11000001";    --SBCI:4
    rom_block(7473)   <=B"0000000000000000_00000010_11000001";    --SBCI:4
    rom_block(7474)   <=B"0000000000000000_00000010_11000001";    --SBCI:4
    rom_block(7475)   <=B"0000000000000000_00000010_11000001";    --SBCI:4
    rom_block(7476)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7477)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7478)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7479)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7480)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7481)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7482)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7483)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7484)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7485)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7486)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7487)   <="00000000000000000000000000000000";    --TBD2:7
    
    rom_block(7488)   <="00000000000000000100000000000100";    --NOP:0
    rom_block(7489)   <="00000000000000000100000000000100";    --NOP:0
    rom_block(7490)   <="00000000000000000100000000000100";    --NOP:0
    rom_block(7491)   <="00000000000000000100000000000100";    --NOP:0
    rom_block(7492)   <="00000000000000000001010000001000";    --NOP:1
    rom_block(7493)   <="00000000000000000001010000001000";    --NOP:1
    rom_block(7494)   <="00000000000000000001010000001000";    --NOP:1
    rom_block(7495)   <="00000000000000000001010000001000";    --NOP:1
    rom_block(7496)   <="00000000000000000000000000000000";    --NOP:2
    rom_block(7497)   <="00000000000000000000000000000000";    --NOP:2
    rom_block(7498)   <="00000000000000000000000000000000";    --NOP:2
    rom_block(7499)   <="00000000000000000000000000000000";    --NOP:2
    rom_block(7500)   <="00000000000000000000000000000000";    --NOP:3
    rom_block(7501)   <="00000000000000000000000000000000";    --NOP:3
    rom_block(7502)   <="00000000000000000000000000000000";    --NOP:3
    rom_block(7503)   <="00000000000000000000000000000000";    --NOP:3
    rom_block(7504)   <="00000000000000000000000000000000";    --NOP:4
    rom_block(7505)   <="00000000000000000000000000000000";    --NOP:4
    rom_block(7506)   <="00000000000000000000000000000000";    --NOP:4
    rom_block(7507)   <="00000000000000000000000000000000";    --NOP:4
    rom_block(7508)   <="00000000000000000000000000000000";    --NOP:5
    rom_block(7509)   <="00000000000000000000000000000000";    --NOP:5
    rom_block(7510)   <="00000000000000000000000000000000";    --NOP:5
    rom_block(7511)   <="00000000000000000000000000000000";    --NOP:5
    rom_block(7512)   <="00000000000000000000000000000000";    --NOP:6
    rom_block(7513)   <="00000000000000000000000000000000";    --NOP:6
    rom_block(7514)   <="00000000000000000000000000000000";    --NOP:6
    rom_block(7515)   <="00000000000000000000000000000000";    --NOP:6
    rom_block(7516)   <="00000000000000000000000000000000";    --NOP:7
    rom_block(7517)   <="00000000000000000000000000000000";    --NOP:7
    rom_block(7518)   <="00000000000000000000000000000000";    --NOP:7
    rom_block(7519)   <="00000000000000000000000000000000";    --NOP:7
    rom_block(7520)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7521)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7522)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7523)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7524)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7525)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7526)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7527)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7528)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7529)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7530)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7531)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7532)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7533)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7534)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7535)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7536)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7537)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7538)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7539)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7540)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7541)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7542)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7543)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7544)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7545)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7546)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7547)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7548)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7549)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7550)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7551)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7552)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7553)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7554)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7555)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7556)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7557)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7558)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7559)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7560)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7561)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7562)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7563)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7564)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7565)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7566)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7567)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7568)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7569)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7570)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7571)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7572)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7573)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7574)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7575)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7576)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7577)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7578)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7579)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7580)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7581)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7582)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7583)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7584)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7585)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7586)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7587)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7588)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7589)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7590)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7591)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7592)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7593)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7594)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7595)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7596)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7597)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7598)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7599)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7600)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7601)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7602)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7603)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7604)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7605)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7606)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7607)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7608)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7609)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7610)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7611)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7612)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7613)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7614)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7615)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7616)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7617)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7618)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7619)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7620)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7621)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7622)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7623)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7624)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7625)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7626)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7627)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7628)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7629)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7630)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7631)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7632)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7633)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7634)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7635)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7636)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7637)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7638)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7639)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7640)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7641)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7642)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7643)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7644)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7645)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7646)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7647)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7648)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7649)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7650)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7651)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7652)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7653)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7654)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7655)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7656)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7657)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7658)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7659)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7660)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7661)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7662)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7663)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7664)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7665)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7666)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7667)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7668)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7669)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7670)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7671)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7672)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7673)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7674)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7675)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7676)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7677)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7678)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7679)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7680)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7681)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7682)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7683)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7684)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7685)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7686)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7687)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7688)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7689)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7690)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7691)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7692)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7693)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7694)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7695)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7696)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7697)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7698)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7699)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7700)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7701)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7702)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7703)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7704)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7705)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7706)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7707)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7708)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7709)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7710)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7711)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7712)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7713)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7714)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7715)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7716)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7717)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7718)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7719)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7720)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7721)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7722)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7723)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7724)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7725)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7726)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7727)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7728)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7729)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7730)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7731)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7732)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7733)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7734)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7735)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7736)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7737)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7738)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7739)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7740)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7741)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7742)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7743)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7744)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7745)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7746)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7747)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7748)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7749)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7750)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7751)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7752)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7753)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7754)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7755)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7756)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7757)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7758)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7759)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7760)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7761)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7762)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7763)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7764)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7765)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7766)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7767)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7768)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7769)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7770)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7771)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7772)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7773)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7774)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7775)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7776)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7777)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7778)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7779)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7780)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7781)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7782)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7783)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7784)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7785)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7786)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7787)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7788)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7789)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7790)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7791)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7792)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7793)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7794)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7795)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7796)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7797)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7798)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7799)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7800)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7801)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7802)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7803)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7804)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7805)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7806)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7807)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7808)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7809)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7810)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7811)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7812)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7813)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7814)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7815)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7816)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7817)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7818)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7819)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7820)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7821)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7822)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7823)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7824)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7825)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7826)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7827)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7828)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7829)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7830)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7831)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7832)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7833)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7834)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7835)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7836)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7837)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7838)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7839)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7840)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7841)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7842)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7843)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7844)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7845)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7846)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7847)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7848)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7849)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7850)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7851)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7852)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7853)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7854)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7855)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7856)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7857)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7858)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7859)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7860)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7861)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7862)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7863)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7864)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7865)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7866)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7867)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7868)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7869)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7870)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7871)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7872)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7873)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7874)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7875)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7876)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7877)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7878)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7879)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7880)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7881)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7882)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7883)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7884)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7885)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7886)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7887)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7888)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7889)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7890)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7891)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7892)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7893)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7894)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7895)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7896)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7897)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7898)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7899)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7900)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7901)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7902)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7903)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7904)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7905)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7906)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7907)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7908)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7909)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7910)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7911)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7912)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7913)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7914)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7915)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7916)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7917)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7918)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7919)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7920)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7921)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7922)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7923)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7924)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7925)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7926)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7927)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7928)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7929)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7930)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7931)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7932)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7933)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7934)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7935)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7936)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7937)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7938)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7939)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(7940)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7941)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7942)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7943)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(7944)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7945)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7946)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7947)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(7948)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7949)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7950)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7951)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(7952)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7953)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7954)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7955)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(7956)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7957)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7958)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7959)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(7960)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7961)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7962)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7963)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(7964)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7965)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7966)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7967)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(7968)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7969)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7970)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7971)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(7972)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7973)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7974)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7975)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(7976)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7977)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7978)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7979)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(7980)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7981)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7982)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7983)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(7984)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7985)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7986)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7987)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(7988)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7989)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7990)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7991)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(7992)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7993)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7994)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7995)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(7996)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7997)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7998)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(7999)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(8000)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8001)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8002)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8003)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8004)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8005)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8006)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8007)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8008)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8009)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8010)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8011)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8012)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8013)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8014)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8015)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8016)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8017)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8018)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8019)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8020)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8021)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8022)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8023)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8024)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8025)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8026)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8027)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8028)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(8029)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(8030)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(8031)   <="00000000000000000000000000000000";    --TBD:7
    
    -- xx/xx/xx/xx/xx/xx/xx/xx
    -- xx/xx/xx/ IOUT / IIN / YOUT / YIN / XOUT 
    -- HLT / MEMADDRIN / RAMIN / RAMOUT / INSTOUT / INSTIN / AIN / AOUT 
    -- SUMOUT / SUBTRACT / XIN / OUTREGIN / COUNTEN (PC++) / COUNTOUT (PC) / JUMP(set PC) / FI   
    --LDI Immediate (FB)
    rom_block(8032)   <=B"00000000_00000000_01000000_00000100";    --LDII:0             -step 0
    rom_block(8033)   <="00000000000000000100000000000100";    --LDII:0
    rom_block(8034)   <="00000000000000000100000000000100";    --LDII:0
    rom_block(8035)   <="00000000000000000100000000000100";    --LDII:0
    rom_block(8036)   <="00000000000000000001010000001000";    --LDII:1             -step 1
    rom_block(8037)   <="00000000000000000001010000001000";    --LDII:1
    rom_block(8038)   <="00000000000000000001010000001000";    --LDII:1
    rom_block(8039)   <="00000000000000000001010000001000";    --LDII:1
    rom_block(8040)   <=B"0000000000000000_0100000000000100";    --LDII:2             -step 2                 
    rom_block(8041)   <=B"0000000000000000_0100000000000100";    --LDII:2
    rom_block(8042)   <=B"0000000000000000_0100000000000100";    --LDII:2
    rom_block(8043)   <=B"0000000000000000_0100000000000100";    --LDII:2
    rom_block(8044)   <=B"0000000000001000_0001000000001000";    --LDII:3
    rom_block(8045)   <=B"0000000000001000_0001000000001000";    --LDII:3
    rom_block(8046)   <=B"0000000000001000_0001000000001000";    --LDII:3
    rom_block(8047)   <=B"0000000000001000_0001000000001000";    --LDII:3
    rom_block(8048)   <="00000000000000000000000000000100";    --LDII:4
    rom_block(8049)   <="00000000000000000000000000000100";    --LDII:4
    rom_block(8050)   <="00000000000000000000000000000100";    --LDII:4
    rom_block(8051)   <="00000000000000000000000000000100";    --LDII:4
    rom_block(8052)   <="00000000000000000000000000000000";    --LDII:5
    rom_block(8053)   <="00000000000000000000000000000000";    --LDII:5
    rom_block(8054)   <="00000000000000000000000000000000";    --LDII:5
    rom_block(8055)   <="00000000000000000000000000000000";    --LDII:5
    rom_block(8056)   <="00000000000000000000000000000000";    --LDII:6
    rom_block(8057)   <="00000000000000000000000000000000";    --LDII:6
    rom_block(8058)   <="00000000000000000000000000000000";    --LDII:6
    rom_block(8059)   <="00000000000000000000000000000000";    --LDII:6
    rom_block(8060)   <="00000000000000000000000000000000";    --LDII:7
    rom_block(8061)   <="00000000000000000000000000000000";    --LDII:7
    rom_block(8062)   <="00000000000000000000000000000000";    --LDII:7
    rom_block(8063)   <="00000000000000000000000000000000";    --LDII:7
    
    rom_block(8064)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8065)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8066)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8067)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8068)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8069)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8070)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8071)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8072)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8073)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8074)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8075)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8076)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8077)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8078)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8079)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8080)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8081)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8082)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8083)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8084)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8085)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8086)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8087)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8088)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8089)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8090)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8091)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8092)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(8093)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(8094)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(8095)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(8096)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(8097)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(8098)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(8099)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(8100)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(8101)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(8102)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(8103)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(8104)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(8105)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(8106)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(8107)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(8108)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(8109)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(8110)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(8111)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(8112)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(8113)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(8114)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(8115)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(8116)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(8117)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(8118)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(8119)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(8120)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(8121)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(8122)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(8123)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(8124)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(8125)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(8126)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(8127)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(8128)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8129)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8130)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8131)   <="00000000000000000100000000000100";    --TBD:0
    rom_block(8132)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8133)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8134)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8135)   <="00000000000000000001010000001000";    --TBD:1
    rom_block(8136)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8137)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8138)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8139)   <="00000000000000000000000000000000";    --TBD:2
    rom_block(8140)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8141)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8142)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8143)   <="00000000000000000000000000000000";    --TBD:3
    rom_block(8144)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8145)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8146)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8147)   <="00000000000000000000000000000000";    --TBD:4
    rom_block(8148)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8149)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8150)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8151)   <="00000000000000000000000000000000";    --TBD:5
    rom_block(8152)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8153)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8154)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8155)   <="00000000000000000000000000000000";    --TBD:6
    rom_block(8156)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(8157)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(8158)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(8159)   <="00000000000000000000000000000000";    --TBD:7
    rom_block(8160)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(8161)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(8162)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(8163)   <="00000000000000000100000000000100";    --TBD2:0
    rom_block(8164)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(8165)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(8166)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(8167)   <="00000000000000000001010000001000";    --TBD2:1
    rom_block(8168)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(8169)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(8170)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(8171)   <="00000000000000000000000000000000";    --TBD2:2
    rom_block(8172)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(8173)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(8174)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(8175)   <="00000000000000000000000000000000";    --TBD2:3
    rom_block(8176)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(8177)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(8178)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(8179)   <="00000000000000000000000000000000";    --TBD2:4
    rom_block(8180)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(8181)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(8182)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(8183)   <="00000000000000000000000000000000";    --TBD2:5
    rom_block(8184)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(8185)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(8186)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(8187)   <="00000000000000000000000000000000";    --TBD2:6
    rom_block(8188)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(8189)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(8190)   <="00000000000000000000000000000000";    --TBD2:7
    rom_block(8191)   <="00000000000000000000000000000000";    --TBD2:7
    
   -- IOUT / IIN / YOUT / YIN / XOUT / HLT / MEMADDRIN / RAMIN / RAMOUT / INSTOUT / INSTIN / AIN / AOUT / SUMOUT / SUBTRACT / XIN / OUTREGIN / COUNTEN (PC++) / COUNTOUT (PC) / JUMP(set PC) / FI
   PROCESS (sys_clk_i, inst, step, flags)
    
   BEGIN
         --addr<=to_integer(shift_left(unsigned(resize(unsigned(inst),8)),4) + unsigned(step));         --IIII0SSS
         --addr <= to_integer(unsigned(inst) & '0' & unsigned(step));
         
         --IIIIIIIISSSFF   Instruction Step Flag
         addr <= to_integer(unsigned(inst) & unsigned(step) & unsigned(flags(1 downto 0)));     --1 carry, 0 zero
         
         q_I_OUT_t                  <= rom_block(addr)(20);
         q_I_IN_t                   <= rom_block(addr)(19);
         q_Y_OUT_t                  <= rom_block(addr)(18);
         q_Y_IN_t                   <= rom_block(addr)(17);
         q_X_OUT_t                  <= rom_block(addr)(16);
         q_HALT_t                   <= rom_block(addr)(15);
         q_MEM_ADDR_IN_t            <= rom_block(addr)(14);
         q_RAM_IN_t                 <= rom_block(addr)(13);
         q_RAM_OUT_t                <= rom_block(addr)(12);
         q_INST_OUT_t               <= rom_block(addr)(11);
         q_INST_IN_t                <= rom_block(addr)(10);
         q_A_IN_t                   <= rom_block(addr)(9);
         q_A_OUT_t                  <= rom_block(addr)(8);
         q_SUM_OUT_t                <= rom_block(addr)(7);
         q_SUBTRACT_t               <= rom_block(addr)(6);
         q_X_IN_t                   <= rom_block(addr)(5);
         q_OUTREG_IN_t              <= rom_block(addr)(4);
         q_COUNTER_ENABLE_t         <= rom_block(addr)(3);
         q_COUNTER_OUT_t            <= rom_block(addr)(2);
         q_JUMP_t                   <= rom_block(addr)(1);
         q_FI_t                     <= rom_block(addr)(0);
    
   END PROCESS;
   
    q_CONTROL16        <= rom_block(addr);
    --q_CurrentADDR      <= std_logic_vector(to_unsigned(addr,9));
    q_CurrentADDR      <= std_logic_vector(to_unsigned(addr,13));
    
    q_I_OUT             <= q_I_OUT_t;
    q_I_IN              <= q_I_IN_t;
    q_Y_OUT             <= q_Y_OUT_t;
    q_Y_IN              <= q_Y_IN_t;
    q_X_OUT             <= q_X_OUT_t; 
    q_HALT              <= q_HALT_t;
    q_MEM_ADDR_IN       <= q_MEM_ADDR_IN_t;
    q_RAM_IN            <= q_RAM_IN_t;
    q_RAM_OUT           <= q_RAM_OUT_t;
    q_INST_OUT          <= q_INST_OUT_t;
    q_INST_IN           <= q_INST_IN_t;
    q_A_IN              <= q_A_IN_t;
    q_A_OUT             <= q_A_OUT_t;
    q_SUM_OUT           <= q_SUM_OUT_t;
    q_SUBTRACT          <= q_SUBTRACT_t;
    q_X_IN              <= q_X_IN_t;
    q_OUTREG_IN         <= q_OUTREG_IN_t;
    q_COUNTER_ENABLE    <= q_COUNTER_ENABLE_t;
    q_COUNTER_OUT       <= q_COUNTER_OUT_t;
    q_JUMP              <= q_JUMP_t;
    q_FI                <= q_FI_t;

end Behavioral;
