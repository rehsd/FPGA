library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

entity BusData is
    Port ( 
        d_in_A                      : IN std_logic_vector (15 downto 0);
        d_in_X                      : IN std_logic_vector (15 downto 0);
        d_in_Y                      : IN std_logic_vector (15 downto 0);
        d_in_I                      : IN std_logic_vector (15 downto 0);
        d_in_SUM                    : IN std_logic_vector (15 downto 0);
        d_in_COUNTER                : IN std_logic_vector (15 downto 0);
        d_in_MEM_ADDR               : IN std_logic_vector (15 downto 0);
        d_in_MEM                    : IN std_logic_vector (15 downto 0);
        d_in_INST                   : IN std_logic_vector (15 downto 0);
        load_enable_A               : IN std_logic;
        load_enable_X               : IN std_logic;
        load_enable_Y               : IN std_logic;
        load_enable_I               : IN std_logic;
        load_enable_SUM             : IN std_logic;
        load_enable_COUNTER         : IN std_logic;
        load_enable_MEM_ADDR        : IN std_logic;
        load_enable_MEM             : IN std_logic;
        load_enable_INST            : IN std_logic;
        load_enable_JMP             : IN std_logic;
        clr                         : IN std_logic;
        sys_clk_i                   : IN std_logic;
        q_out                       : OUT std_logic_vector (15 downto 0)  := "0000000000000000"
    );
end BusData;
    
architecture Behavioral of BusData is
    signal tempOut: std_logic_vector (15 downto 0) := "0000000000000000";
begin
    process(d_in_A, d_in_X, d_in_Y, d_in_I, d_in_SUM, d_in_COUNTER, d_in_MEM_ADDR, d_in_MEM, d_in_INST, load_enable_A, load_enable_X, load_enable_Y, load_enable_I, 
        load_enable_SUM, load_enable_COUNTER, load_enable_MEM_ADDR, load_enable_MEM, load_enable_INST, clr, sys_clk_i, load_enable_JMP)
    begin 
        if(clr='1') then
            tempOut <="0000000000000000";
        else --if(rising_edge(sys_clk_i)) then
            if (load_enable_COUNTER = '1') then
                tempOut <= d_in_COUNTER;
            elsif(load_enable_MEM = '1') then 
                tempOut <=d_in_MEM;
            elsif load_enable_A = '1' then
                tempOut <= d_in_A ;
            elsif load_enable_X = '1' then
                tempOut <= d_in_X;
            elsif load_enable_Y = '1' then
                tempOut <= d_in_Y;
            elsif load_enable_I = '1' then
                tempOut <= d_in_I;
            elsif load_enable_SUM = '1' then
                tempOut <= d_in_SUM ;
            elsif load_enable_MEM_ADDR  = '1' then
                tempOut <= d_in_MEM_ADDR;
            elsif load_enable_INST  = '1' then
                tempOut <= d_in_INST  ;
            elsif load_enable_JMP = '1' then
                tempOut <= d_in_MEM;
            else
                tempOut <= tempOut;     
            end if;
        end if;
    end process;
    q_out<=tempOut;
end Behavioral;
