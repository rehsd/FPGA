
`timescale 1 ns / 1 ps

	module rehsd_gfx_writer #
	(
		// Users to add parameters here

		// User parameters ends
		
		//parameter  C_M00_AXI_START_DATA_VALUE	= 32'hFF00FFFF,
		//parameter  C_M00_AXI_TARGET_SLAVE_BASE_ADDR	= 32'h30900000,
		parameter integer C_M00_AXI_ADDR_WIDTH	= 32,
		parameter integer C_M00_AXI_DATA_WIDTH	= 32,
		parameter integer C_M00_AXI_TRANSACTIONS_NUM	= 1
	)
	(
		// Users to add ports here
        input wire [31:0] addr_to_write,
        input wire [31:0] color_to_write,
		// User ports ends

		// Ports of Axi Master Bus Interface M00_AXI
		input wire  m00_axi_init_axi_txn,
		output wire  m00_axi_error,
		output wire  m00_axi_txn_done,
		input wire  m00_axi_aclk,
		input wire  m00_axi_aresetn,
		output wire [C_M00_AXI_ADDR_WIDTH-1 : 0] m00_axi_awaddr,
		output wire [2 : 0] m00_axi_awprot,
		output wire  m00_axi_awvalid,
		input wire  m00_axi_awready,
		output wire [C_M00_AXI_DATA_WIDTH-1 : 0] m00_axi_wdata,
		output wire [C_M00_AXI_DATA_WIDTH/8-1 : 0] m00_axi_wstrb,
		output wire  m00_axi_wvalid,
		input wire  m00_axi_wready,
		input wire [1 : 0] m00_axi_bresp,
		input wire  m00_axi_bvalid,
		output wire  m00_axi_bready,
		output wire [C_M00_AXI_ADDR_WIDTH-1 : 0] m00_axi_araddr,
		output wire [2 : 0] m00_axi_arprot,
		output wire  m00_axi_arvalid,
		input wire  m00_axi_arready,
		input wire [C_M00_AXI_DATA_WIDTH-1 : 0] m00_axi_rdata,
		input wire [1 : 0] m00_axi_rresp,
		input wire  m00_axi_rvalid,
		output wire  m00_axi_rready
	);
	
	//use registers so that if addr/color change mid-cycle, they remain a set
	reg [31:0] addr_reg;
    reg [31:0] color_reg;
    reg m00_axi_init_axi_txn_prev;
    
    always @(posedge m00_axi_aclk) begin
        if (!m00_axi_init_axi_txn_prev && m00_axi_init_axi_txn) begin
            addr_reg  <= addr_to_write;
            color_reg <= color_to_write;
        end
        m00_axi_init_axi_txn_prev <= m00_axi_init_axi_txn; // Store previous state
    end 

// Instantiation of Axi Bus Interface M00_AXI
	rehsd_gfx_writer_master_lite_v1_0_M00_AXI # ( 
		//.C_M_START_DATA_VALUE(32'hFFFFFFFF),
		//.C_M_TARGET_SLAVE_BASE_ADDR(32'h30900000),
		.C_M_AXI_ADDR_WIDTH(C_M00_AXI_ADDR_WIDTH),
		.C_M_AXI_DATA_WIDTH(C_M00_AXI_DATA_WIDTH),
		.C_M_TRANSACTIONS_NUM(C_M00_AXI_TRANSACTIONS_NUM)
	) rehsd_gfx_writer_master_lite_v1_0_M00_AXI_inst (
		.addr_to_write(addr_reg),
		.color_to_write(color_reg),
		.INIT_AXI_TXN(m00_axi_init_axi_txn),
		.ERROR(m00_axi_error),
		.TXN_DONE(m00_axi_txn_done),
		.M_AXI_ACLK(m00_axi_aclk),
		.M_AXI_ARESETN(m00_axi_aresetn),
		.M_AXI_AWADDR(m00_axi_awaddr),
		.M_AXI_AWPROT(m00_axi_awprot),
		.M_AXI_AWVALID(m00_axi_awvalid),
		.M_AXI_AWREADY(m00_axi_awready),
		.M_AXI_WDATA(m00_axi_wdata),
		.M_AXI_WSTRB(m00_axi_wstrb),
		.M_AXI_WVALID(m00_axi_wvalid),
		.M_AXI_WREADY(m00_axi_wready),
		.M_AXI_BRESP(m00_axi_bresp),
		.M_AXI_BVALID(m00_axi_bvalid),
		.M_AXI_BREADY(m00_axi_bready),
		.M_AXI_ARADDR(m00_axi_araddr),
		.M_AXI_ARPROT(m00_axi_arprot),
		.M_AXI_ARVALID(m00_axi_arvalid),
		.M_AXI_ARREADY(m00_axi_arready),
		.M_AXI_RDATA(m00_axi_rdata),
		.M_AXI_RRESP(m00_axi_rresp),
		.M_AXI_RVALID(m00_axi_rvalid),
		.M_AXI_RREADY(m00_axi_rready)
	);

	// Add user logic here
    
    
	// User logic ends

	endmodule